module top (
    // 16MHz clock
    input CLK,

    // USB pull-up resistor
    output USBPU,

    // R1, G1, B1
    output PIN_1,
    output PIN_2,
    output PIN_3,
    output PIN_4,
    output PIN_5

);

    // drive USB pull-up resistor to '0' to disable USB
    assign USBPU = 0;

    wire clk_10mhz;
    assign PIN_1 = red;
    assign PIN_2 = green;
    assign PIN_3 = blue;
    assign PIN_4 = h_sync;
    assign PIN_5 = v_sync;

    reg [8:0] h_counter;
    reg [0:0] h_sync;

    reg [9:0] v_counter;
    reg [0:0] v_sync;

    reg [0:0] red;
    reg [0:0] green;
    reg [0:0] blue;

    // Create a 10MHz clock.
    // http://martin.hinner.info/vga/timing.html
    // 40 MHz = 800x600@60Hz
    // 10 MHz = 200x150
    SB_PLL40_CORE #(
      .DIVR(0),
      .DIVF(9),
      .DIVQ(4),
      .FILTER_RANGE(3'b001),
      .FEEDBACK_PATH("SIMPLE"),
      .DELAY_ADJUSTMENT_MODE_FEEDBACK("FIXED"),
      .FDA_FEEDBACK(4'b0000),
      .DELAY_ADJUSTMENT_MODE_RELATIVE("FIXED"),
      .FDA_RELATIVE(4'b0000),
      .SHIFTREG_DIV_MODE(2'b00),
      .PLLOUT_SELECT("GENCLK"),
      .ENABLE_ICEGATE(1'b0)
    ) pll (
      .REFERENCECLK(CLK),
      .PLLOUTCORE(clk_10mhz),
      .RESETB(1),
      .BYPASS(0)
    );

    reg [2:0] memory_array [0:30000];

    // Zero out display.
    initial begin
      $readmemb("memory_array.mem", memory_array);

      memory_array[0] <= 3'b111;
      memory_array[1] <= 3'b111;
      memory_array[2] <= 3'b111;
      memory_array[3] <= 3'b111;
      memory_array[4] <= 3'b111;
      memory_array[5] <= 3'b111;
      memory_array[6] <= 3'b111;
      memory_array[7] <= 3'b111;
      memory_array[8] <= 3'b101;
      memory_array[9] <= 3'b101;
      memory_array[10] <= 3'b000;
      memory_array[11] <= 3'b101;
      memory_array[12] <= 3'b101;
      memory_array[13] <= 3'b101;
      memory_array[14] <= 3'b101;
      memory_array[15] <= 3'b101;
      memory_array[16] <= 3'b101;
      memory_array[17] <= 3'b000;
      memory_array[18] <= 3'b101;
      memory_array[19] <= 3'b101;
      memory_array[20] <= 3'b000;
      memory_array[21] <= 3'b101;
      memory_array[22] <= 3'b101;
      memory_array[23] <= 3'b101;
      memory_array[24] <= 3'b101;
      memory_array[25] <= 3'b101;
      memory_array[26] <= 3'b101;
      memory_array[27] <= 3'b000;
      memory_array[28] <= 3'b101;
      memory_array[29] <= 3'b101;
      memory_array[30] <= 3'b000;
      memory_array[31] <= 3'b101;
      memory_array[32] <= 3'b101;
      memory_array[33] <= 3'b101;
      memory_array[34] <= 3'b101;
      memory_array[35] <= 3'b101;
      memory_array[36] <= 3'b101;
      memory_array[37] <= 3'b000;
      memory_array[38] <= 3'b101;
      memory_array[39] <= 3'b101;
      memory_array[40] <= 3'b000;
      memory_array[41] <= 3'b101;
      memory_array[42] <= 3'b101;
      memory_array[43] <= 3'b101;
      memory_array[44] <= 3'b101;
      memory_array[45] <= 3'b101;
      memory_array[46] <= 3'b101;
      memory_array[47] <= 3'b000;
      memory_array[48] <= 3'b101;
      memory_array[49] <= 3'b101;
      memory_array[50] <= 3'b000;
      memory_array[51] <= 3'b101;
      memory_array[52] <= 3'b101;
      memory_array[53] <= 3'b101;
      memory_array[54] <= 3'b101;
      memory_array[55] <= 3'b101;
      memory_array[56] <= 3'b101;
      memory_array[57] <= 3'b000;
      memory_array[58] <= 3'b101;
      memory_array[59] <= 3'b101;
      memory_array[60] <= 3'b000;
      memory_array[61] <= 3'b101;
      memory_array[62] <= 3'b101;
      memory_array[63] <= 3'b101;
      memory_array[64] <= 3'b101;
      memory_array[65] <= 3'b101;
      memory_array[66] <= 3'b101;
      memory_array[67] <= 3'b000;
      memory_array[68] <= 3'b101;
      memory_array[69] <= 3'b101;
      memory_array[70] <= 3'b000;
      memory_array[71] <= 3'b101;
      memory_array[72] <= 3'b101;
      memory_array[73] <= 3'b101;
      memory_array[74] <= 3'b101;
      memory_array[75] <= 3'b101;
      memory_array[76] <= 3'b101;
      memory_array[77] <= 3'b000;
      memory_array[78] <= 3'b101;
      memory_array[79] <= 3'b101;
      memory_array[80] <= 3'b000;
      memory_array[81] <= 3'b101;
      memory_array[82] <= 3'b101;
      memory_array[83] <= 3'b101;
      memory_array[84] <= 3'b101;
      memory_array[85] <= 3'b101;
      memory_array[86] <= 3'b101;
      memory_array[87] <= 3'b000;
      memory_array[88] <= 3'b101;
      memory_array[89] <= 3'b101;
      memory_array[90] <= 3'b000;
      memory_array[91] <= 3'b101;
      memory_array[92] <= 3'b101;
      memory_array[93] <= 3'b101;
      memory_array[94] <= 3'b000;
      memory_array[95] <= 3'b111;
      memory_array[96] <= 3'b111;
      memory_array[97] <= 3'b111;
      memory_array[98] <= 3'b111;
      memory_array[99] <= 3'b000;
      memory_array[100] <= 3'b000;
      memory_array[101] <= 3'b111;
      memory_array[102] <= 3'b111;
      memory_array[103] <= 3'b111;
      memory_array[104] <= 3'b111;
      memory_array[105] <= 3'b000;
      memory_array[106] <= 3'b101;
      memory_array[107] <= 3'b101;
      memory_array[108] <= 3'b101;
      memory_array[109] <= 3'b110;
      memory_array[110] <= 3'b101;
      memory_array[111] <= 3'b101;
      memory_array[112] <= 3'b101;
      memory_array[113] <= 3'b101;
      memory_array[114] <= 3'b101;
      memory_array[115] <= 3'b101;
      memory_array[116] <= 3'b101;
      memory_array[117] <= 3'b101;
      memory_array[118] <= 3'b101;
      memory_array[119] <= 3'b110;
      memory_array[120] <= 3'b101;
      memory_array[121] <= 3'b101;
      memory_array[122] <= 3'b101;
      memory_array[123] <= 3'b101;
      memory_array[124] <= 3'b101;
      memory_array[125] <= 3'b101;
      memory_array[126] <= 3'b101;
      memory_array[127] <= 3'b101;
      memory_array[128] <= 3'b101;
      memory_array[129] <= 3'b110;
      memory_array[130] <= 3'b101;
      memory_array[131] <= 3'b101;
      memory_array[132] <= 3'b101;
      memory_array[133] <= 3'b101;
      memory_array[134] <= 3'b101;
      memory_array[135] <= 3'b101;
      memory_array[136] <= 3'b101;
      memory_array[137] <= 3'b101;
      memory_array[138] <= 3'b101;
      memory_array[139] <= 3'b110;
      memory_array[140] <= 3'b101;
      memory_array[141] <= 3'b101;
      memory_array[142] <= 3'b101;
      memory_array[143] <= 3'b101;
      memory_array[144] <= 3'b101;
      memory_array[145] <= 3'b101;
      memory_array[146] <= 3'b101;
      memory_array[147] <= 3'b101;
      memory_array[148] <= 3'b101;
      memory_array[149] <= 3'b110;
      memory_array[150] <= 3'b101;
      memory_array[151] <= 3'b101;
      memory_array[152] <= 3'b101;
      memory_array[153] <= 3'b101;
      memory_array[154] <= 3'b101;
      memory_array[155] <= 3'b101;
      memory_array[156] <= 3'b101;
      memory_array[157] <= 3'b101;
      memory_array[158] <= 3'b101;
      memory_array[159] <= 3'b110;
      memory_array[160] <= 3'b101;
      memory_array[161] <= 3'b101;
      memory_array[162] <= 3'b101;
      memory_array[163] <= 3'b101;
      memory_array[164] <= 3'b101;
      memory_array[165] <= 3'b101;
      memory_array[166] <= 3'b101;
      memory_array[167] <= 3'b101;
      memory_array[168] <= 3'b101;
      memory_array[169] <= 3'b110;
      memory_array[170] <= 3'b101;
      memory_array[171] <= 3'b101;
      memory_array[172] <= 3'b101;
      memory_array[173] <= 3'b101;
      memory_array[174] <= 3'b101;
      memory_array[175] <= 3'b101;
      memory_array[176] <= 3'b101;
      memory_array[177] <= 3'b101;
      memory_array[178] <= 3'b101;
      memory_array[179] <= 3'b110;
      memory_array[180] <= 3'b101;
      memory_array[181] <= 3'b101;
      memory_array[182] <= 3'b101;
      memory_array[183] <= 3'b101;
      memory_array[184] <= 3'b101;
      memory_array[185] <= 3'b101;
      memory_array[186] <= 3'b101;
      memory_array[187] <= 3'b101;
      memory_array[188] <= 3'b101;
      memory_array[189] <= 3'b110;
      memory_array[190] <= 3'b101;
      memory_array[191] <= 3'b101;
      memory_array[192] <= 3'b111;
      memory_array[193] <= 3'b111;
      memory_array[194] <= 3'b111;
      memory_array[195] <= 3'b111;
      memory_array[196] <= 3'b111;
      memory_array[197] <= 3'b111;
      memory_array[198] <= 3'b111;
      memory_array[199] <= 3'b111;
      memory_array[200] <= 3'b111;
      memory_array[201] <= 3'b111;
      memory_array[202] <= 3'b111;
      memory_array[203] <= 3'b111;
      memory_array[204] <= 3'b111;
      memory_array[205] <= 3'b111;
      memory_array[206] <= 3'b111;
      memory_array[207] <= 3'b111;
      memory_array[208] <= 3'b101;
      memory_array[209] <= 3'b101;
      memory_array[210] <= 3'b110;
      memory_array[211] <= 3'b101;
      memory_array[212] <= 3'b101;
      memory_array[213] <= 3'b101;
      memory_array[214] <= 3'b101;
      memory_array[215] <= 3'b101;
      memory_array[216] <= 3'b101;
      memory_array[217] <= 3'b110;
      memory_array[218] <= 3'b101;
      memory_array[219] <= 3'b101;
      memory_array[220] <= 3'b110;
      memory_array[221] <= 3'b101;
      memory_array[222] <= 3'b101;
      memory_array[223] <= 3'b101;
      memory_array[224] <= 3'b101;
      memory_array[225] <= 3'b101;
      memory_array[226] <= 3'b101;
      memory_array[227] <= 3'b110;
      memory_array[228] <= 3'b101;
      memory_array[229] <= 3'b101;
      memory_array[230] <= 3'b110;
      memory_array[231] <= 3'b101;
      memory_array[232] <= 3'b101;
      memory_array[233] <= 3'b101;
      memory_array[234] <= 3'b101;
      memory_array[235] <= 3'b101;
      memory_array[236] <= 3'b101;
      memory_array[237] <= 3'b110;
      memory_array[238] <= 3'b101;
      memory_array[239] <= 3'b101;
      memory_array[240] <= 3'b110;
      memory_array[241] <= 3'b101;
      memory_array[242] <= 3'b101;
      memory_array[243] <= 3'b101;
      memory_array[244] <= 3'b101;
      memory_array[245] <= 3'b101;
      memory_array[246] <= 3'b101;
      memory_array[247] <= 3'b110;
      memory_array[248] <= 3'b101;
      memory_array[249] <= 3'b101;
      memory_array[250] <= 3'b110;
      memory_array[251] <= 3'b101;
      memory_array[252] <= 3'b101;
      memory_array[253] <= 3'b101;
      memory_array[254] <= 3'b101;
      memory_array[255] <= 3'b101;
      memory_array[256] <= 3'b101;
      memory_array[257] <= 3'b110;
      memory_array[258] <= 3'b101;
      memory_array[259] <= 3'b101;
      memory_array[260] <= 3'b110;
      memory_array[261] <= 3'b101;
      memory_array[262] <= 3'b101;
      memory_array[263] <= 3'b101;
      memory_array[264] <= 3'b101;
      memory_array[265] <= 3'b101;
      memory_array[266] <= 3'b101;
      memory_array[267] <= 3'b110;
      memory_array[268] <= 3'b101;
      memory_array[269] <= 3'b101;
      memory_array[270] <= 3'b110;
      memory_array[271] <= 3'b101;
      memory_array[272] <= 3'b101;
      memory_array[273] <= 3'b101;
      memory_array[274] <= 3'b101;
      memory_array[275] <= 3'b101;
      memory_array[276] <= 3'b101;
      memory_array[277] <= 3'b110;
      memory_array[278] <= 3'b101;
      memory_array[279] <= 3'b101;
      memory_array[280] <= 3'b110;
      memory_array[281] <= 3'b101;
      memory_array[282] <= 3'b101;
      memory_array[283] <= 3'b101;
      memory_array[284] <= 3'b101;
      memory_array[285] <= 3'b101;
      memory_array[286] <= 3'b101;
      memory_array[287] <= 3'b110;
      memory_array[288] <= 3'b101;
      memory_array[289] <= 3'b101;
      memory_array[290] <= 3'b110;
      memory_array[291] <= 3'b101;
      memory_array[292] <= 3'b101;
      memory_array[293] <= 3'b101;
      memory_array[294] <= 3'b000;
      memory_array[295] <= 3'b101;
      memory_array[296] <= 3'b111;
      memory_array[297] <= 3'b111;
      memory_array[298] <= 3'b111;
      memory_array[299] <= 3'b000;
      memory_array[300] <= 3'b000;
      memory_array[301] <= 3'b111;
      memory_array[302] <= 3'b111;
      memory_array[303] <= 3'b111;
      memory_array[304] <= 3'b101;
      memory_array[305] <= 3'b000;
      memory_array[306] <= 3'b101;
      memory_array[307] <= 3'b101;
      memory_array[308] <= 3'b101;
      memory_array[309] <= 3'b000;
      memory_array[310] <= 3'b101;
      memory_array[311] <= 3'b101;
      memory_array[312] <= 3'b110;
      memory_array[313] <= 3'b101;
      memory_array[314] <= 3'b101;
      memory_array[315] <= 3'b101;
      memory_array[316] <= 3'b101;
      memory_array[317] <= 3'b101;
      memory_array[318] <= 3'b101;
      memory_array[319] <= 3'b000;
      memory_array[320] <= 3'b101;
      memory_array[321] <= 3'b101;
      memory_array[322] <= 3'b110;
      memory_array[323] <= 3'b101;
      memory_array[324] <= 3'b101;
      memory_array[325] <= 3'b101;
      memory_array[326] <= 3'b101;
      memory_array[327] <= 3'b101;
      memory_array[328] <= 3'b101;
      memory_array[329] <= 3'b000;
      memory_array[330] <= 3'b101;
      memory_array[331] <= 3'b101;
      memory_array[332] <= 3'b110;
      memory_array[333] <= 3'b101;
      memory_array[334] <= 3'b101;
      memory_array[335] <= 3'b101;
      memory_array[336] <= 3'b101;
      memory_array[337] <= 3'b101;
      memory_array[338] <= 3'b101;
      memory_array[339] <= 3'b000;
      memory_array[340] <= 3'b101;
      memory_array[341] <= 3'b101;
      memory_array[342] <= 3'b110;
      memory_array[343] <= 3'b101;
      memory_array[344] <= 3'b101;
      memory_array[345] <= 3'b101;
      memory_array[346] <= 3'b101;
      memory_array[347] <= 3'b101;
      memory_array[348] <= 3'b101;
      memory_array[349] <= 3'b000;
      memory_array[350] <= 3'b101;
      memory_array[351] <= 3'b101;
      memory_array[352] <= 3'b110;
      memory_array[353] <= 3'b101;
      memory_array[354] <= 3'b101;
      memory_array[355] <= 3'b101;
      memory_array[356] <= 3'b101;
      memory_array[357] <= 3'b101;
      memory_array[358] <= 3'b101;
      memory_array[359] <= 3'b000;
      memory_array[360] <= 3'b101;
      memory_array[361] <= 3'b101;
      memory_array[362] <= 3'b110;
      memory_array[363] <= 3'b101;
      memory_array[364] <= 3'b101;
      memory_array[365] <= 3'b101;
      memory_array[366] <= 3'b101;
      memory_array[367] <= 3'b101;
      memory_array[368] <= 3'b101;
      memory_array[369] <= 3'b000;
      memory_array[370] <= 3'b101;
      memory_array[371] <= 3'b101;
      memory_array[372] <= 3'b110;
      memory_array[373] <= 3'b101;
      memory_array[374] <= 3'b101;
      memory_array[375] <= 3'b101;
      memory_array[376] <= 3'b101;
      memory_array[377] <= 3'b101;
      memory_array[378] <= 3'b101;
      memory_array[379] <= 3'b000;
      memory_array[380] <= 3'b101;
      memory_array[381] <= 3'b101;
      memory_array[382] <= 3'b110;
      memory_array[383] <= 3'b101;
      memory_array[384] <= 3'b101;
      memory_array[385] <= 3'b101;
      memory_array[386] <= 3'b101;
      memory_array[387] <= 3'b101;
      memory_array[388] <= 3'b101;
      memory_array[389] <= 3'b000;
      memory_array[390] <= 3'b101;
      memory_array[391] <= 3'b101;
      memory_array[392] <= 3'b111;
      memory_array[393] <= 3'b111;
      memory_array[394] <= 3'b111;
      memory_array[395] <= 3'b111;
      memory_array[396] <= 3'b111;
      memory_array[397] <= 3'b111;
      memory_array[398] <= 3'b111;
      memory_array[399] <= 3'b111;
      memory_array[400] <= 3'b111;
      memory_array[401] <= 3'b111;
      memory_array[402] <= 3'b111;
      memory_array[403] <= 3'b101;
      memory_array[404] <= 3'b101;
      memory_array[405] <= 3'b111;
      memory_array[406] <= 3'b111;
      memory_array[407] <= 3'b111;
      memory_array[408] <= 3'b101;
      memory_array[409] <= 3'b101;
      memory_array[410] <= 3'b110;
      memory_array[411] <= 3'b110;
      memory_array[412] <= 3'b101;
      memory_array[413] <= 3'b101;
      memory_array[414] <= 3'b101;
      memory_array[415] <= 3'b101;
      memory_array[416] <= 3'b110;
      memory_array[417] <= 3'b110;
      memory_array[418] <= 3'b101;
      memory_array[419] <= 3'b101;
      memory_array[420] <= 3'b110;
      memory_array[421] <= 3'b110;
      memory_array[422] <= 3'b101;
      memory_array[423] <= 3'b101;
      memory_array[424] <= 3'b101;
      memory_array[425] <= 3'b101;
      memory_array[426] <= 3'b110;
      memory_array[427] <= 3'b110;
      memory_array[428] <= 3'b101;
      memory_array[429] <= 3'b101;
      memory_array[430] <= 3'b110;
      memory_array[431] <= 3'b110;
      memory_array[432] <= 3'b101;
      memory_array[433] <= 3'b101;
      memory_array[434] <= 3'b101;
      memory_array[435] <= 3'b101;
      memory_array[436] <= 3'b110;
      memory_array[437] <= 3'b110;
      memory_array[438] <= 3'b101;
      memory_array[439] <= 3'b101;
      memory_array[440] <= 3'b110;
      memory_array[441] <= 3'b110;
      memory_array[442] <= 3'b101;
      memory_array[443] <= 3'b101;
      memory_array[444] <= 3'b101;
      memory_array[445] <= 3'b101;
      memory_array[446] <= 3'b110;
      memory_array[447] <= 3'b110;
      memory_array[448] <= 3'b101;
      memory_array[449] <= 3'b101;
      memory_array[450] <= 3'b110;
      memory_array[451] <= 3'b110;
      memory_array[452] <= 3'b101;
      memory_array[453] <= 3'b101;
      memory_array[454] <= 3'b101;
      memory_array[455] <= 3'b101;
      memory_array[456] <= 3'b110;
      memory_array[457] <= 3'b110;
      memory_array[458] <= 3'b101;
      memory_array[459] <= 3'b101;
      memory_array[460] <= 3'b110;
      memory_array[461] <= 3'b110;
      memory_array[462] <= 3'b101;
      memory_array[463] <= 3'b101;
      memory_array[464] <= 3'b101;
      memory_array[465] <= 3'b101;
      memory_array[466] <= 3'b110;
      memory_array[467] <= 3'b110;
      memory_array[468] <= 3'b101;
      memory_array[469] <= 3'b101;
      memory_array[470] <= 3'b110;
      memory_array[471] <= 3'b110;
      memory_array[472] <= 3'b101;
      memory_array[473] <= 3'b101;
      memory_array[474] <= 3'b101;
      memory_array[475] <= 3'b101;
      memory_array[476] <= 3'b110;
      memory_array[477] <= 3'b110;
      memory_array[478] <= 3'b101;
      memory_array[479] <= 3'b101;
      memory_array[480] <= 3'b110;
      memory_array[481] <= 3'b110;
      memory_array[482] <= 3'b101;
      memory_array[483] <= 3'b101;
      memory_array[484] <= 3'b101;
      memory_array[485] <= 3'b101;
      memory_array[486] <= 3'b110;
      memory_array[487] <= 3'b110;
      memory_array[488] <= 3'b101;
      memory_array[489] <= 3'b101;
      memory_array[490] <= 3'b110;
      memory_array[491] <= 3'b110;
      memory_array[492] <= 3'b101;
      memory_array[493] <= 3'b101;
      memory_array[494] <= 3'b000;
      memory_array[495] <= 3'b101;
      memory_array[496] <= 3'b111;
      memory_array[497] <= 3'b111;
      memory_array[498] <= 3'b111;
      memory_array[499] <= 3'b000;
      memory_array[500] <= 3'b000;
      memory_array[501] <= 3'b111;
      memory_array[502] <= 3'b111;
      memory_array[503] <= 3'b111;
      memory_array[504] <= 3'b101;
      memory_array[505] <= 3'b000;
      memory_array[506] <= 3'b101;
      memory_array[507] <= 3'b110;
      memory_array[508] <= 3'b000;
      memory_array[509] <= 3'b000;
      memory_array[510] <= 3'b101;
      memory_array[511] <= 3'b101;
      memory_array[512] <= 3'b110;
      memory_array[513] <= 3'b000;
      memory_array[514] <= 3'b101;
      memory_array[515] <= 3'b101;
      memory_array[516] <= 3'b101;
      memory_array[517] <= 3'b110;
      memory_array[518] <= 3'b000;
      memory_array[519] <= 3'b000;
      memory_array[520] <= 3'b101;
      memory_array[521] <= 3'b101;
      memory_array[522] <= 3'b110;
      memory_array[523] <= 3'b000;
      memory_array[524] <= 3'b101;
      memory_array[525] <= 3'b101;
      memory_array[526] <= 3'b101;
      memory_array[527] <= 3'b110;
      memory_array[528] <= 3'b000;
      memory_array[529] <= 3'b000;
      memory_array[530] <= 3'b101;
      memory_array[531] <= 3'b101;
      memory_array[532] <= 3'b110;
      memory_array[533] <= 3'b000;
      memory_array[534] <= 3'b101;
      memory_array[535] <= 3'b101;
      memory_array[536] <= 3'b101;
      memory_array[537] <= 3'b110;
      memory_array[538] <= 3'b000;
      memory_array[539] <= 3'b000;
      memory_array[540] <= 3'b101;
      memory_array[541] <= 3'b101;
      memory_array[542] <= 3'b110;
      memory_array[543] <= 3'b000;
      memory_array[544] <= 3'b101;
      memory_array[545] <= 3'b101;
      memory_array[546] <= 3'b101;
      memory_array[547] <= 3'b110;
      memory_array[548] <= 3'b000;
      memory_array[549] <= 3'b000;
      memory_array[550] <= 3'b101;
      memory_array[551] <= 3'b101;
      memory_array[552] <= 3'b110;
      memory_array[553] <= 3'b000;
      memory_array[554] <= 3'b101;
      memory_array[555] <= 3'b101;
      memory_array[556] <= 3'b101;
      memory_array[557] <= 3'b110;
      memory_array[558] <= 3'b000;
      memory_array[559] <= 3'b000;
      memory_array[560] <= 3'b101;
      memory_array[561] <= 3'b101;
      memory_array[562] <= 3'b110;
      memory_array[563] <= 3'b000;
      memory_array[564] <= 3'b101;
      memory_array[565] <= 3'b101;
      memory_array[566] <= 3'b101;
      memory_array[567] <= 3'b110;
      memory_array[568] <= 3'b000;
      memory_array[569] <= 3'b000;
      memory_array[570] <= 3'b101;
      memory_array[571] <= 3'b101;
      memory_array[572] <= 3'b110;
      memory_array[573] <= 3'b000;
      memory_array[574] <= 3'b101;
      memory_array[575] <= 3'b101;
      memory_array[576] <= 3'b101;
      memory_array[577] <= 3'b110;
      memory_array[578] <= 3'b000;
      memory_array[579] <= 3'b000;
      memory_array[580] <= 3'b101;
      memory_array[581] <= 3'b101;
      memory_array[582] <= 3'b110;
      memory_array[583] <= 3'b000;
      memory_array[584] <= 3'b101;
      memory_array[585] <= 3'b101;
      memory_array[586] <= 3'b101;
      memory_array[587] <= 3'b110;
      memory_array[588] <= 3'b000;
      memory_array[589] <= 3'b000;
      memory_array[590] <= 3'b101;
      memory_array[591] <= 3'b101;
      memory_array[592] <= 3'b111;
      memory_array[593] <= 3'b111;
      memory_array[594] <= 3'b111;
      memory_array[595] <= 3'b101;
      memory_array[596] <= 3'b101;
      memory_array[597] <= 3'b111;
      memory_array[598] <= 3'b111;
      memory_array[599] <= 3'b111;
      memory_array[600] <= 3'b111;
      memory_array[601] <= 3'b111;
      memory_array[602] <= 3'b111;
      memory_array[603] <= 3'b101;
      memory_array[604] <= 3'b101;
      memory_array[605] <= 3'b111;
      memory_array[606] <= 3'b111;
      memory_array[607] <= 3'b111;
      memory_array[608] <= 3'b101;
      memory_array[609] <= 3'b101;
      memory_array[610] <= 3'b000;
      memory_array[611] <= 3'b000;
      memory_array[612] <= 3'b101;
      memory_array[613] <= 3'b101;
      memory_array[614] <= 3'b101;
      memory_array[615] <= 3'b101;
      memory_array[616] <= 3'b000;
      memory_array[617] <= 3'b000;
      memory_array[618] <= 3'b101;
      memory_array[619] <= 3'b101;
      memory_array[620] <= 3'b000;
      memory_array[621] <= 3'b000;
      memory_array[622] <= 3'b101;
      memory_array[623] <= 3'b101;
      memory_array[624] <= 3'b101;
      memory_array[625] <= 3'b101;
      memory_array[626] <= 3'b000;
      memory_array[627] <= 3'b000;
      memory_array[628] <= 3'b101;
      memory_array[629] <= 3'b101;
      memory_array[630] <= 3'b000;
      memory_array[631] <= 3'b000;
      memory_array[632] <= 3'b101;
      memory_array[633] <= 3'b101;
      memory_array[634] <= 3'b101;
      memory_array[635] <= 3'b101;
      memory_array[636] <= 3'b000;
      memory_array[637] <= 3'b000;
      memory_array[638] <= 3'b101;
      memory_array[639] <= 3'b101;
      memory_array[640] <= 3'b000;
      memory_array[641] <= 3'b000;
      memory_array[642] <= 3'b101;
      memory_array[643] <= 3'b101;
      memory_array[644] <= 3'b101;
      memory_array[645] <= 3'b101;
      memory_array[646] <= 3'b000;
      memory_array[647] <= 3'b000;
      memory_array[648] <= 3'b101;
      memory_array[649] <= 3'b101;
      memory_array[650] <= 3'b000;
      memory_array[651] <= 3'b000;
      memory_array[652] <= 3'b101;
      memory_array[653] <= 3'b101;
      memory_array[654] <= 3'b101;
      memory_array[655] <= 3'b101;
      memory_array[656] <= 3'b000;
      memory_array[657] <= 3'b000;
      memory_array[658] <= 3'b101;
      memory_array[659] <= 3'b101;
      memory_array[660] <= 3'b000;
      memory_array[661] <= 3'b000;
      memory_array[662] <= 3'b101;
      memory_array[663] <= 3'b101;
      memory_array[664] <= 3'b101;
      memory_array[665] <= 3'b101;
      memory_array[666] <= 3'b000;
      memory_array[667] <= 3'b000;
      memory_array[668] <= 3'b101;
      memory_array[669] <= 3'b101;
      memory_array[670] <= 3'b000;
      memory_array[671] <= 3'b000;
      memory_array[672] <= 3'b101;
      memory_array[673] <= 3'b101;
      memory_array[674] <= 3'b101;
      memory_array[675] <= 3'b101;
      memory_array[676] <= 3'b000;
      memory_array[677] <= 3'b000;
      memory_array[678] <= 3'b101;
      memory_array[679] <= 3'b101;
      memory_array[680] <= 3'b000;
      memory_array[681] <= 3'b000;
      memory_array[682] <= 3'b101;
      memory_array[683] <= 3'b101;
      memory_array[684] <= 3'b101;
      memory_array[685] <= 3'b101;
      memory_array[686] <= 3'b000;
      memory_array[687] <= 3'b000;
      memory_array[688] <= 3'b101;
      memory_array[689] <= 3'b101;
      memory_array[690] <= 3'b000;
      memory_array[691] <= 3'b000;
      memory_array[692] <= 3'b101;
      memory_array[693] <= 3'b101;
      memory_array[694] <= 3'b000;
      memory_array[695] <= 3'b101;
      memory_array[696] <= 3'b111;
      memory_array[697] <= 3'b111;
      memory_array[698] <= 3'b111;
      memory_array[699] <= 3'b000;
      memory_array[700] <= 3'b000;
      memory_array[701] <= 3'b111;
      memory_array[702] <= 3'b111;
      memory_array[703] <= 3'b111;
      memory_array[704] <= 3'b101;
      memory_array[705] <= 3'b000;
      memory_array[706] <= 3'b101;
      memory_array[707] <= 3'b000;
      memory_array[708] <= 3'b110;
      memory_array[709] <= 3'b110;
      memory_array[710] <= 3'b101;
      memory_array[711] <= 3'b101;
      memory_array[712] <= 3'b000;
      memory_array[713] <= 3'b110;
      memory_array[714] <= 3'b101;
      memory_array[715] <= 3'b101;
      memory_array[716] <= 3'b101;
      memory_array[717] <= 3'b000;
      memory_array[718] <= 3'b110;
      memory_array[719] <= 3'b110;
      memory_array[720] <= 3'b101;
      memory_array[721] <= 3'b101;
      memory_array[722] <= 3'b000;
      memory_array[723] <= 3'b110;
      memory_array[724] <= 3'b101;
      memory_array[725] <= 3'b101;
      memory_array[726] <= 3'b101;
      memory_array[727] <= 3'b000;
      memory_array[728] <= 3'b110;
      memory_array[729] <= 3'b110;
      memory_array[730] <= 3'b101;
      memory_array[731] <= 3'b101;
      memory_array[732] <= 3'b000;
      memory_array[733] <= 3'b110;
      memory_array[734] <= 3'b101;
      memory_array[735] <= 3'b101;
      memory_array[736] <= 3'b101;
      memory_array[737] <= 3'b000;
      memory_array[738] <= 3'b110;
      memory_array[739] <= 3'b110;
      memory_array[740] <= 3'b101;
      memory_array[741] <= 3'b101;
      memory_array[742] <= 3'b000;
      memory_array[743] <= 3'b110;
      memory_array[744] <= 3'b101;
      memory_array[745] <= 3'b101;
      memory_array[746] <= 3'b101;
      memory_array[747] <= 3'b000;
      memory_array[748] <= 3'b110;
      memory_array[749] <= 3'b110;
      memory_array[750] <= 3'b101;
      memory_array[751] <= 3'b101;
      memory_array[752] <= 3'b000;
      memory_array[753] <= 3'b110;
      memory_array[754] <= 3'b101;
      memory_array[755] <= 3'b101;
      memory_array[756] <= 3'b101;
      memory_array[757] <= 3'b000;
      memory_array[758] <= 3'b110;
      memory_array[759] <= 3'b110;
      memory_array[760] <= 3'b101;
      memory_array[761] <= 3'b101;
      memory_array[762] <= 3'b000;
      memory_array[763] <= 3'b110;
      memory_array[764] <= 3'b101;
      memory_array[765] <= 3'b101;
      memory_array[766] <= 3'b101;
      memory_array[767] <= 3'b000;
      memory_array[768] <= 3'b110;
      memory_array[769] <= 3'b110;
      memory_array[770] <= 3'b101;
      memory_array[771] <= 3'b101;
      memory_array[772] <= 3'b000;
      memory_array[773] <= 3'b110;
      memory_array[774] <= 3'b101;
      memory_array[775] <= 3'b101;
      memory_array[776] <= 3'b101;
      memory_array[777] <= 3'b000;
      memory_array[778] <= 3'b110;
      memory_array[779] <= 3'b110;
      memory_array[780] <= 3'b101;
      memory_array[781] <= 3'b101;
      memory_array[782] <= 3'b000;
      memory_array[783] <= 3'b110;
      memory_array[784] <= 3'b101;
      memory_array[785] <= 3'b101;
      memory_array[786] <= 3'b101;
      memory_array[787] <= 3'b000;
      memory_array[788] <= 3'b110;
      memory_array[789] <= 3'b110;
      memory_array[790] <= 3'b101;
      memory_array[791] <= 3'b101;
      memory_array[792] <= 3'b111;
      memory_array[793] <= 3'b111;
      memory_array[794] <= 3'b111;
      memory_array[795] <= 3'b101;
      memory_array[796] <= 3'b101;
      memory_array[797] <= 3'b111;
      memory_array[798] <= 3'b111;
      memory_array[799] <= 3'b111;
      memory_array[800] <= 3'b111;
      memory_array[801] <= 3'b101;
      memory_array[802] <= 3'b101;
      memory_array[803] <= 3'b111;
      memory_array[804] <= 3'b111;
      memory_array[805] <= 3'b101;
      memory_array[806] <= 3'b101;
      memory_array[807] <= 3'b111;
      memory_array[808] <= 3'b101;
      memory_array[809] <= 3'b101;
      memory_array[810] <= 3'b000;
      memory_array[811] <= 3'b101;
      memory_array[812] <= 3'b111;
      memory_array[813] <= 3'b111;
      memory_array[814] <= 3'b111;
      memory_array[815] <= 3'b111;
      memory_array[816] <= 3'b101;
      memory_array[817] <= 3'b000;
      memory_array[818] <= 3'b101;
      memory_array[819] <= 3'b101;
      memory_array[820] <= 3'b000;
      memory_array[821] <= 3'b101;
      memory_array[822] <= 3'b111;
      memory_array[823] <= 3'b111;
      memory_array[824] <= 3'b111;
      memory_array[825] <= 3'b111;
      memory_array[826] <= 3'b101;
      memory_array[827] <= 3'b000;
      memory_array[828] <= 3'b101;
      memory_array[829] <= 3'b101;
      memory_array[830] <= 3'b000;
      memory_array[831] <= 3'b101;
      memory_array[832] <= 3'b111;
      memory_array[833] <= 3'b111;
      memory_array[834] <= 3'b111;
      memory_array[835] <= 3'b111;
      memory_array[836] <= 3'b101;
      memory_array[837] <= 3'b000;
      memory_array[838] <= 3'b101;
      memory_array[839] <= 3'b101;
      memory_array[840] <= 3'b000;
      memory_array[841] <= 3'b101;
      memory_array[842] <= 3'b111;
      memory_array[843] <= 3'b111;
      memory_array[844] <= 3'b111;
      memory_array[845] <= 3'b111;
      memory_array[846] <= 3'b101;
      memory_array[847] <= 3'b000;
      memory_array[848] <= 3'b101;
      memory_array[849] <= 3'b101;
      memory_array[850] <= 3'b000;
      memory_array[851] <= 3'b101;
      memory_array[852] <= 3'b111;
      memory_array[853] <= 3'b111;
      memory_array[854] <= 3'b111;
      memory_array[855] <= 3'b111;
      memory_array[856] <= 3'b101;
      memory_array[857] <= 3'b000;
      memory_array[858] <= 3'b101;
      memory_array[859] <= 3'b101;
      memory_array[860] <= 3'b000;
      memory_array[861] <= 3'b101;
      memory_array[862] <= 3'b111;
      memory_array[863] <= 3'b111;
      memory_array[864] <= 3'b111;
      memory_array[865] <= 3'b111;
      memory_array[866] <= 3'b101;
      memory_array[867] <= 3'b000;
      memory_array[868] <= 3'b101;
      memory_array[869] <= 3'b101;
      memory_array[870] <= 3'b000;
      memory_array[871] <= 3'b101;
      memory_array[872] <= 3'b111;
      memory_array[873] <= 3'b111;
      memory_array[874] <= 3'b111;
      memory_array[875] <= 3'b111;
      memory_array[876] <= 3'b101;
      memory_array[877] <= 3'b000;
      memory_array[878] <= 3'b101;
      memory_array[879] <= 3'b101;
      memory_array[880] <= 3'b000;
      memory_array[881] <= 3'b101;
      memory_array[882] <= 3'b111;
      memory_array[883] <= 3'b111;
      memory_array[884] <= 3'b111;
      memory_array[885] <= 3'b111;
      memory_array[886] <= 3'b101;
      memory_array[887] <= 3'b000;
      memory_array[888] <= 3'b101;
      memory_array[889] <= 3'b101;
      memory_array[890] <= 3'b000;
      memory_array[891] <= 3'b101;
      memory_array[892] <= 3'b111;
      memory_array[893] <= 3'b111;
      memory_array[894] <= 3'b101;
      memory_array[895] <= 3'b111;
      memory_array[896] <= 3'b111;
      memory_array[897] <= 3'b111;
      memory_array[898] <= 3'b111;
      memory_array[899] <= 3'b101;
      memory_array[900] <= 3'b000;
      memory_array[901] <= 3'b111;
      memory_array[902] <= 3'b111;
      memory_array[903] <= 3'b111;
      memory_array[904] <= 3'b111;
      memory_array[905] <= 3'b101;
      memory_array[906] <= 3'b111;
      memory_array[907] <= 3'b111;
      memory_array[908] <= 3'b101;
      memory_array[909] <= 3'b110;
      memory_array[910] <= 3'b101;
      memory_array[911] <= 3'b101;
      memory_array[912] <= 3'b111;
      memory_array[913] <= 3'b101;
      memory_array[914] <= 3'b111;
      memory_array[915] <= 3'b111;
      memory_array[916] <= 3'b111;
      memory_array[917] <= 3'b111;
      memory_array[918] <= 3'b101;
      memory_array[919] <= 3'b110;
      memory_array[920] <= 3'b101;
      memory_array[921] <= 3'b101;
      memory_array[922] <= 3'b111;
      memory_array[923] <= 3'b101;
      memory_array[924] <= 3'b111;
      memory_array[925] <= 3'b111;
      memory_array[926] <= 3'b111;
      memory_array[927] <= 3'b111;
      memory_array[928] <= 3'b101;
      memory_array[929] <= 3'b110;
      memory_array[930] <= 3'b101;
      memory_array[931] <= 3'b101;
      memory_array[932] <= 3'b111;
      memory_array[933] <= 3'b101;
      memory_array[934] <= 3'b111;
      memory_array[935] <= 3'b111;
      memory_array[936] <= 3'b111;
      memory_array[937] <= 3'b111;
      memory_array[938] <= 3'b101;
      memory_array[939] <= 3'b110;
      memory_array[940] <= 3'b101;
      memory_array[941] <= 3'b101;
      memory_array[942] <= 3'b111;
      memory_array[943] <= 3'b101;
      memory_array[944] <= 3'b111;
      memory_array[945] <= 3'b111;
      memory_array[946] <= 3'b111;
      memory_array[947] <= 3'b111;
      memory_array[948] <= 3'b101;
      memory_array[949] <= 3'b110;
      memory_array[950] <= 3'b101;
      memory_array[951] <= 3'b101;
      memory_array[952] <= 3'b111;
      memory_array[953] <= 3'b101;
      memory_array[954] <= 3'b111;
      memory_array[955] <= 3'b111;
      memory_array[956] <= 3'b111;
      memory_array[957] <= 3'b111;
      memory_array[958] <= 3'b101;
      memory_array[959] <= 3'b110;
      memory_array[960] <= 3'b101;
      memory_array[961] <= 3'b101;
      memory_array[962] <= 3'b111;
      memory_array[963] <= 3'b101;
      memory_array[964] <= 3'b111;
      memory_array[965] <= 3'b111;
      memory_array[966] <= 3'b111;
      memory_array[967] <= 3'b111;
      memory_array[968] <= 3'b101;
      memory_array[969] <= 3'b110;
      memory_array[970] <= 3'b101;
      memory_array[971] <= 3'b101;
      memory_array[972] <= 3'b111;
      memory_array[973] <= 3'b101;
      memory_array[974] <= 3'b111;
      memory_array[975] <= 3'b111;
      memory_array[976] <= 3'b111;
      memory_array[977] <= 3'b111;
      memory_array[978] <= 3'b101;
      memory_array[979] <= 3'b110;
      memory_array[980] <= 3'b101;
      memory_array[981] <= 3'b101;
      memory_array[982] <= 3'b111;
      memory_array[983] <= 3'b101;
      memory_array[984] <= 3'b111;
      memory_array[985] <= 3'b111;
      memory_array[986] <= 3'b111;
      memory_array[987] <= 3'b111;
      memory_array[988] <= 3'b101;
      memory_array[989] <= 3'b110;
      memory_array[990] <= 3'b101;
      memory_array[991] <= 3'b101;
      memory_array[992] <= 3'b111;
      memory_array[993] <= 3'b101;
      memory_array[994] <= 3'b101;
      memory_array[995] <= 3'b111;
      memory_array[996] <= 3'b111;
      memory_array[997] <= 3'b101;
      memory_array[998] <= 3'b101;
      memory_array[999] <= 3'b111;
      memory_array[1000] <= 3'b111;
      memory_array[1001] <= 3'b101;
      memory_array[1002] <= 3'b101;
      memory_array[1003] <= 3'b111;
      memory_array[1004] <= 3'b111;
      memory_array[1005] <= 3'b101;
      memory_array[1006] <= 3'b101;
      memory_array[1007] <= 3'b111;
      memory_array[1008] <= 3'b101;
      memory_array[1009] <= 3'b101;
      memory_array[1010] <= 3'b000;
      memory_array[1011] <= 3'b101;
      memory_array[1012] <= 3'b111;
      memory_array[1013] <= 3'b111;
      memory_array[1014] <= 3'b111;
      memory_array[1015] <= 3'b111;
      memory_array[1016] <= 3'b101;
      memory_array[1017] <= 3'b000;
      memory_array[1018] <= 3'b101;
      memory_array[1019] <= 3'b101;
      memory_array[1020] <= 3'b000;
      memory_array[1021] <= 3'b101;
      memory_array[1022] <= 3'b111;
      memory_array[1023] <= 3'b111;
      memory_array[1024] <= 3'b111;
      memory_array[1025] <= 3'b111;
      memory_array[1026] <= 3'b101;
      memory_array[1027] <= 3'b000;
      memory_array[1028] <= 3'b101;
      memory_array[1029] <= 3'b101;
      memory_array[1030] <= 3'b000;
      memory_array[1031] <= 3'b101;
      memory_array[1032] <= 3'b111;
      memory_array[1033] <= 3'b111;
      memory_array[1034] <= 3'b111;
      memory_array[1035] <= 3'b111;
      memory_array[1036] <= 3'b101;
      memory_array[1037] <= 3'b000;
      memory_array[1038] <= 3'b101;
      memory_array[1039] <= 3'b101;
      memory_array[1040] <= 3'b000;
      memory_array[1041] <= 3'b101;
      memory_array[1042] <= 3'b111;
      memory_array[1043] <= 3'b111;
      memory_array[1044] <= 3'b111;
      memory_array[1045] <= 3'b111;
      memory_array[1046] <= 3'b101;
      memory_array[1047] <= 3'b000;
      memory_array[1048] <= 3'b101;
      memory_array[1049] <= 3'b101;
      memory_array[1050] <= 3'b000;
      memory_array[1051] <= 3'b101;
      memory_array[1052] <= 3'b111;
      memory_array[1053] <= 3'b111;
      memory_array[1054] <= 3'b111;
      memory_array[1055] <= 3'b111;
      memory_array[1056] <= 3'b101;
      memory_array[1057] <= 3'b000;
      memory_array[1058] <= 3'b101;
      memory_array[1059] <= 3'b101;
      memory_array[1060] <= 3'b000;
      memory_array[1061] <= 3'b101;
      memory_array[1062] <= 3'b111;
      memory_array[1063] <= 3'b111;
      memory_array[1064] <= 3'b111;
      memory_array[1065] <= 3'b111;
      memory_array[1066] <= 3'b101;
      memory_array[1067] <= 3'b000;
      memory_array[1068] <= 3'b101;
      memory_array[1069] <= 3'b101;
      memory_array[1070] <= 3'b000;
      memory_array[1071] <= 3'b101;
      memory_array[1072] <= 3'b111;
      memory_array[1073] <= 3'b111;
      memory_array[1074] <= 3'b111;
      memory_array[1075] <= 3'b111;
      memory_array[1076] <= 3'b101;
      memory_array[1077] <= 3'b000;
      memory_array[1078] <= 3'b101;
      memory_array[1079] <= 3'b101;
      memory_array[1080] <= 3'b000;
      memory_array[1081] <= 3'b101;
      memory_array[1082] <= 3'b111;
      memory_array[1083] <= 3'b111;
      memory_array[1084] <= 3'b111;
      memory_array[1085] <= 3'b111;
      memory_array[1086] <= 3'b101;
      memory_array[1087] <= 3'b000;
      memory_array[1088] <= 3'b101;
      memory_array[1089] <= 3'b101;
      memory_array[1090] <= 3'b000;
      memory_array[1091] <= 3'b101;
      memory_array[1092] <= 3'b111;
      memory_array[1093] <= 3'b111;
      memory_array[1094] <= 3'b101;
      memory_array[1095] <= 3'b111;
      memory_array[1096] <= 3'b111;
      memory_array[1097] <= 3'b111;
      memory_array[1098] <= 3'b111;
      memory_array[1099] <= 3'b101;
      memory_array[1100] <= 3'b000;
      memory_array[1101] <= 3'b111;
      memory_array[1102] <= 3'b111;
      memory_array[1103] <= 3'b111;
      memory_array[1104] <= 3'b111;
      memory_array[1105] <= 3'b101;
      memory_array[1106] <= 3'b111;
      memory_array[1107] <= 3'b111;
      memory_array[1108] <= 3'b101;
      memory_array[1109] <= 3'b110;
      memory_array[1110] <= 3'b101;
      memory_array[1111] <= 3'b101;
      memory_array[1112] <= 3'b111;
      memory_array[1113] <= 3'b101;
      memory_array[1114] <= 3'b111;
      memory_array[1115] <= 3'b111;
      memory_array[1116] <= 3'b111;
      memory_array[1117] <= 3'b111;
      memory_array[1118] <= 3'b101;
      memory_array[1119] <= 3'b110;
      memory_array[1120] <= 3'b101;
      memory_array[1121] <= 3'b101;
      memory_array[1122] <= 3'b111;
      memory_array[1123] <= 3'b101;
      memory_array[1124] <= 3'b111;
      memory_array[1125] <= 3'b111;
      memory_array[1126] <= 3'b111;
      memory_array[1127] <= 3'b111;
      memory_array[1128] <= 3'b101;
      memory_array[1129] <= 3'b110;
      memory_array[1130] <= 3'b101;
      memory_array[1131] <= 3'b101;
      memory_array[1132] <= 3'b111;
      memory_array[1133] <= 3'b101;
      memory_array[1134] <= 3'b111;
      memory_array[1135] <= 3'b111;
      memory_array[1136] <= 3'b111;
      memory_array[1137] <= 3'b111;
      memory_array[1138] <= 3'b101;
      memory_array[1139] <= 3'b110;
      memory_array[1140] <= 3'b101;
      memory_array[1141] <= 3'b101;
      memory_array[1142] <= 3'b111;
      memory_array[1143] <= 3'b101;
      memory_array[1144] <= 3'b111;
      memory_array[1145] <= 3'b111;
      memory_array[1146] <= 3'b111;
      memory_array[1147] <= 3'b111;
      memory_array[1148] <= 3'b101;
      memory_array[1149] <= 3'b110;
      memory_array[1150] <= 3'b101;
      memory_array[1151] <= 3'b101;
      memory_array[1152] <= 3'b111;
      memory_array[1153] <= 3'b101;
      memory_array[1154] <= 3'b111;
      memory_array[1155] <= 3'b111;
      memory_array[1156] <= 3'b111;
      memory_array[1157] <= 3'b111;
      memory_array[1158] <= 3'b101;
      memory_array[1159] <= 3'b110;
      memory_array[1160] <= 3'b101;
      memory_array[1161] <= 3'b101;
      memory_array[1162] <= 3'b111;
      memory_array[1163] <= 3'b101;
      memory_array[1164] <= 3'b111;
      memory_array[1165] <= 3'b111;
      memory_array[1166] <= 3'b111;
      memory_array[1167] <= 3'b111;
      memory_array[1168] <= 3'b101;
      memory_array[1169] <= 3'b110;
      memory_array[1170] <= 3'b101;
      memory_array[1171] <= 3'b101;
      memory_array[1172] <= 3'b111;
      memory_array[1173] <= 3'b101;
      memory_array[1174] <= 3'b111;
      memory_array[1175] <= 3'b111;
      memory_array[1176] <= 3'b111;
      memory_array[1177] <= 3'b111;
      memory_array[1178] <= 3'b101;
      memory_array[1179] <= 3'b110;
      memory_array[1180] <= 3'b101;
      memory_array[1181] <= 3'b101;
      memory_array[1182] <= 3'b111;
      memory_array[1183] <= 3'b101;
      memory_array[1184] <= 3'b111;
      memory_array[1185] <= 3'b111;
      memory_array[1186] <= 3'b111;
      memory_array[1187] <= 3'b111;
      memory_array[1188] <= 3'b101;
      memory_array[1189] <= 3'b110;
      memory_array[1190] <= 3'b101;
      memory_array[1191] <= 3'b101;
      memory_array[1192] <= 3'b111;
      memory_array[1193] <= 3'b101;
      memory_array[1194] <= 3'b101;
      memory_array[1195] <= 3'b111;
      memory_array[1196] <= 3'b111;
      memory_array[1197] <= 3'b101;
      memory_array[1198] <= 3'b101;
      memory_array[1199] <= 3'b111;
      memory_array[1200] <= 3'b111;
      memory_array[1201] <= 3'b111;
      memory_array[1202] <= 3'b111;
      memory_array[1203] <= 3'b101;
      memory_array[1204] <= 3'b101;
      memory_array[1205] <= 3'b111;
      memory_array[1206] <= 3'b111;
      memory_array[1207] <= 3'b111;
      memory_array[1208] <= 3'b101;
      memory_array[1209] <= 3'b101;
      memory_array[1210] <= 3'b000;
      memory_array[1211] <= 3'b000;
      memory_array[1212] <= 3'b101;
      memory_array[1213] <= 3'b101;
      memory_array[1214] <= 3'b101;
      memory_array[1215] <= 3'b101;
      memory_array[1216] <= 3'b000;
      memory_array[1217] <= 3'b000;
      memory_array[1218] <= 3'b101;
      memory_array[1219] <= 3'b101;
      memory_array[1220] <= 3'b000;
      memory_array[1221] <= 3'b000;
      memory_array[1222] <= 3'b101;
      memory_array[1223] <= 3'b101;
      memory_array[1224] <= 3'b101;
      memory_array[1225] <= 3'b101;
      memory_array[1226] <= 3'b000;
      memory_array[1227] <= 3'b000;
      memory_array[1228] <= 3'b101;
      memory_array[1229] <= 3'b101;
      memory_array[1230] <= 3'b000;
      memory_array[1231] <= 3'b000;
      memory_array[1232] <= 3'b101;
      memory_array[1233] <= 3'b101;
      memory_array[1234] <= 3'b101;
      memory_array[1235] <= 3'b101;
      memory_array[1236] <= 3'b000;
      memory_array[1237] <= 3'b000;
      memory_array[1238] <= 3'b101;
      memory_array[1239] <= 3'b101;
      memory_array[1240] <= 3'b000;
      memory_array[1241] <= 3'b000;
      memory_array[1242] <= 3'b101;
      memory_array[1243] <= 3'b101;
      memory_array[1244] <= 3'b101;
      memory_array[1245] <= 3'b101;
      memory_array[1246] <= 3'b000;
      memory_array[1247] <= 3'b000;
      memory_array[1248] <= 3'b101;
      memory_array[1249] <= 3'b101;
      memory_array[1250] <= 3'b000;
      memory_array[1251] <= 3'b000;
      memory_array[1252] <= 3'b101;
      memory_array[1253] <= 3'b101;
      memory_array[1254] <= 3'b101;
      memory_array[1255] <= 3'b101;
      memory_array[1256] <= 3'b000;
      memory_array[1257] <= 3'b000;
      memory_array[1258] <= 3'b101;
      memory_array[1259] <= 3'b101;
      memory_array[1260] <= 3'b000;
      memory_array[1261] <= 3'b000;
      memory_array[1262] <= 3'b101;
      memory_array[1263] <= 3'b101;
      memory_array[1264] <= 3'b101;
      memory_array[1265] <= 3'b101;
      memory_array[1266] <= 3'b000;
      memory_array[1267] <= 3'b000;
      memory_array[1268] <= 3'b101;
      memory_array[1269] <= 3'b101;
      memory_array[1270] <= 3'b000;
      memory_array[1271] <= 3'b000;
      memory_array[1272] <= 3'b101;
      memory_array[1273] <= 3'b101;
      memory_array[1274] <= 3'b101;
      memory_array[1275] <= 3'b101;
      memory_array[1276] <= 3'b000;
      memory_array[1277] <= 3'b000;
      memory_array[1278] <= 3'b101;
      memory_array[1279] <= 3'b101;
      memory_array[1280] <= 3'b000;
      memory_array[1281] <= 3'b000;
      memory_array[1282] <= 3'b101;
      memory_array[1283] <= 3'b101;
      memory_array[1284] <= 3'b101;
      memory_array[1285] <= 3'b101;
      memory_array[1286] <= 3'b000;
      memory_array[1287] <= 3'b000;
      memory_array[1288] <= 3'b101;
      memory_array[1289] <= 3'b101;
      memory_array[1290] <= 3'b000;
      memory_array[1291] <= 3'b000;
      memory_array[1292] <= 3'b101;
      memory_array[1293] <= 3'b000;
      memory_array[1294] <= 3'b111;
      memory_array[1295] <= 3'b111;
      memory_array[1296] <= 3'b111;
      memory_array[1297] <= 3'b111;
      memory_array[1298] <= 3'b101;
      memory_array[1299] <= 3'b101;
      memory_array[1300] <= 3'b000;
      memory_array[1301] <= 3'b101;
      memory_array[1302] <= 3'b111;
      memory_array[1303] <= 3'b111;
      memory_array[1304] <= 3'b111;
      memory_array[1305] <= 3'b111;
      memory_array[1306] <= 3'b000;
      memory_array[1307] <= 3'b000;
      memory_array[1308] <= 3'b110;
      memory_array[1309] <= 3'b110;
      memory_array[1310] <= 3'b101;
      memory_array[1311] <= 3'b101;
      memory_array[1312] <= 3'b000;
      memory_array[1313] <= 3'b110;
      memory_array[1314] <= 3'b101;
      memory_array[1315] <= 3'b101;
      memory_array[1316] <= 3'b101;
      memory_array[1317] <= 3'b000;
      memory_array[1318] <= 3'b110;
      memory_array[1319] <= 3'b110;
      memory_array[1320] <= 3'b101;
      memory_array[1321] <= 3'b101;
      memory_array[1322] <= 3'b000;
      memory_array[1323] <= 3'b110;
      memory_array[1324] <= 3'b101;
      memory_array[1325] <= 3'b101;
      memory_array[1326] <= 3'b101;
      memory_array[1327] <= 3'b000;
      memory_array[1328] <= 3'b110;
      memory_array[1329] <= 3'b110;
      memory_array[1330] <= 3'b101;
      memory_array[1331] <= 3'b101;
      memory_array[1332] <= 3'b000;
      memory_array[1333] <= 3'b110;
      memory_array[1334] <= 3'b101;
      memory_array[1335] <= 3'b101;
      memory_array[1336] <= 3'b101;
      memory_array[1337] <= 3'b000;
      memory_array[1338] <= 3'b110;
      memory_array[1339] <= 3'b110;
      memory_array[1340] <= 3'b101;
      memory_array[1341] <= 3'b101;
      memory_array[1342] <= 3'b000;
      memory_array[1343] <= 3'b110;
      memory_array[1344] <= 3'b101;
      memory_array[1345] <= 3'b101;
      memory_array[1346] <= 3'b101;
      memory_array[1347] <= 3'b000;
      memory_array[1348] <= 3'b110;
      memory_array[1349] <= 3'b110;
      memory_array[1350] <= 3'b101;
      memory_array[1351] <= 3'b101;
      memory_array[1352] <= 3'b000;
      memory_array[1353] <= 3'b110;
      memory_array[1354] <= 3'b101;
      memory_array[1355] <= 3'b101;
      memory_array[1356] <= 3'b101;
      memory_array[1357] <= 3'b000;
      memory_array[1358] <= 3'b110;
      memory_array[1359] <= 3'b110;
      memory_array[1360] <= 3'b101;
      memory_array[1361] <= 3'b101;
      memory_array[1362] <= 3'b000;
      memory_array[1363] <= 3'b110;
      memory_array[1364] <= 3'b101;
      memory_array[1365] <= 3'b101;
      memory_array[1366] <= 3'b101;
      memory_array[1367] <= 3'b000;
      memory_array[1368] <= 3'b110;
      memory_array[1369] <= 3'b110;
      memory_array[1370] <= 3'b101;
      memory_array[1371] <= 3'b101;
      memory_array[1372] <= 3'b000;
      memory_array[1373] <= 3'b110;
      memory_array[1374] <= 3'b101;
      memory_array[1375] <= 3'b101;
      memory_array[1376] <= 3'b101;
      memory_array[1377] <= 3'b000;
      memory_array[1378] <= 3'b110;
      memory_array[1379] <= 3'b110;
      memory_array[1380] <= 3'b101;
      memory_array[1381] <= 3'b101;
      memory_array[1382] <= 3'b000;
      memory_array[1383] <= 3'b110;
      memory_array[1384] <= 3'b101;
      memory_array[1385] <= 3'b101;
      memory_array[1386] <= 3'b101;
      memory_array[1387] <= 3'b000;
      memory_array[1388] <= 3'b110;
      memory_array[1389] <= 3'b110;
      memory_array[1390] <= 3'b101;
      memory_array[1391] <= 3'b101;
      memory_array[1392] <= 3'b111;
      memory_array[1393] <= 3'b111;
      memory_array[1394] <= 3'b111;
      memory_array[1395] <= 3'b101;
      memory_array[1396] <= 3'b101;
      memory_array[1397] <= 3'b111;
      memory_array[1398] <= 3'b111;
      memory_array[1399] <= 3'b111;
      memory_array[1400] <= 3'b111;
      memory_array[1401] <= 3'b111;
      memory_array[1402] <= 3'b111;
      memory_array[1403] <= 3'b101;
      memory_array[1404] <= 3'b101;
      memory_array[1405] <= 3'b111;
      memory_array[1406] <= 3'b111;
      memory_array[1407] <= 3'b111;
      memory_array[1408] <= 3'b101;
      memory_array[1409] <= 3'b101;
      memory_array[1410] <= 3'b000;
      memory_array[1411] <= 3'b000;
      memory_array[1412] <= 3'b101;
      memory_array[1413] <= 3'b101;
      memory_array[1414] <= 3'b101;
      memory_array[1415] <= 3'b101;
      memory_array[1416] <= 3'b000;
      memory_array[1417] <= 3'b000;
      memory_array[1418] <= 3'b101;
      memory_array[1419] <= 3'b101;
      memory_array[1420] <= 3'b000;
      memory_array[1421] <= 3'b000;
      memory_array[1422] <= 3'b101;
      memory_array[1423] <= 3'b101;
      memory_array[1424] <= 3'b101;
      memory_array[1425] <= 3'b101;
      memory_array[1426] <= 3'b000;
      memory_array[1427] <= 3'b000;
      memory_array[1428] <= 3'b101;
      memory_array[1429] <= 3'b101;
      memory_array[1430] <= 3'b000;
      memory_array[1431] <= 3'b000;
      memory_array[1432] <= 3'b101;
      memory_array[1433] <= 3'b101;
      memory_array[1434] <= 3'b101;
      memory_array[1435] <= 3'b101;
      memory_array[1436] <= 3'b000;
      memory_array[1437] <= 3'b000;
      memory_array[1438] <= 3'b101;
      memory_array[1439] <= 3'b101;
      memory_array[1440] <= 3'b000;
      memory_array[1441] <= 3'b000;
      memory_array[1442] <= 3'b101;
      memory_array[1443] <= 3'b101;
      memory_array[1444] <= 3'b101;
      memory_array[1445] <= 3'b101;
      memory_array[1446] <= 3'b000;
      memory_array[1447] <= 3'b000;
      memory_array[1448] <= 3'b101;
      memory_array[1449] <= 3'b101;
      memory_array[1450] <= 3'b000;
      memory_array[1451] <= 3'b000;
      memory_array[1452] <= 3'b101;
      memory_array[1453] <= 3'b101;
      memory_array[1454] <= 3'b101;
      memory_array[1455] <= 3'b101;
      memory_array[1456] <= 3'b000;
      memory_array[1457] <= 3'b000;
      memory_array[1458] <= 3'b101;
      memory_array[1459] <= 3'b101;
      memory_array[1460] <= 3'b000;
      memory_array[1461] <= 3'b000;
      memory_array[1462] <= 3'b101;
      memory_array[1463] <= 3'b101;
      memory_array[1464] <= 3'b101;
      memory_array[1465] <= 3'b101;
      memory_array[1466] <= 3'b000;
      memory_array[1467] <= 3'b000;
      memory_array[1468] <= 3'b101;
      memory_array[1469] <= 3'b101;
      memory_array[1470] <= 3'b000;
      memory_array[1471] <= 3'b000;
      memory_array[1472] <= 3'b101;
      memory_array[1473] <= 3'b101;
      memory_array[1474] <= 3'b101;
      memory_array[1475] <= 3'b101;
      memory_array[1476] <= 3'b000;
      memory_array[1477] <= 3'b000;
      memory_array[1478] <= 3'b101;
      memory_array[1479] <= 3'b101;
      memory_array[1480] <= 3'b000;
      memory_array[1481] <= 3'b000;
      memory_array[1482] <= 3'b101;
      memory_array[1483] <= 3'b101;
      memory_array[1484] <= 3'b101;
      memory_array[1485] <= 3'b101;
      memory_array[1486] <= 3'b000;
      memory_array[1487] <= 3'b000;
      memory_array[1488] <= 3'b101;
      memory_array[1489] <= 3'b101;
      memory_array[1490] <= 3'b000;
      memory_array[1491] <= 3'b000;
      memory_array[1492] <= 3'b000;
      memory_array[1493] <= 3'b101;
      memory_array[1494] <= 3'b111;
      memory_array[1495] <= 3'b111;
      memory_array[1496] <= 3'b111;
      memory_array[1497] <= 3'b101;
      memory_array[1498] <= 3'b000;
      memory_array[1499] <= 3'b101;
      memory_array[1500] <= 3'b000;
      memory_array[1501] <= 3'b000;
      memory_array[1502] <= 3'b111;
      memory_array[1503] <= 3'b111;
      memory_array[1504] <= 3'b111;
      memory_array[1505] <= 3'b111;
      memory_array[1506] <= 3'b101;
      memory_array[1507] <= 3'b000;
      memory_array[1508] <= 3'b110;
      memory_array[1509] <= 3'b110;
      memory_array[1510] <= 3'b101;
      memory_array[1511] <= 3'b101;
      memory_array[1512] <= 3'b000;
      memory_array[1513] <= 3'b110;
      memory_array[1514] <= 3'b101;
      memory_array[1515] <= 3'b101;
      memory_array[1516] <= 3'b101;
      memory_array[1517] <= 3'b101;
      memory_array[1518] <= 3'b110;
      memory_array[1519] <= 3'b110;
      memory_array[1520] <= 3'b101;
      memory_array[1521] <= 3'b101;
      memory_array[1522] <= 3'b000;
      memory_array[1523] <= 3'b110;
      memory_array[1524] <= 3'b101;
      memory_array[1525] <= 3'b101;
      memory_array[1526] <= 3'b101;
      memory_array[1527] <= 3'b101;
      memory_array[1528] <= 3'b110;
      memory_array[1529] <= 3'b110;
      memory_array[1530] <= 3'b101;
      memory_array[1531] <= 3'b101;
      memory_array[1532] <= 3'b000;
      memory_array[1533] <= 3'b110;
      memory_array[1534] <= 3'b101;
      memory_array[1535] <= 3'b101;
      memory_array[1536] <= 3'b101;
      memory_array[1537] <= 3'b101;
      memory_array[1538] <= 3'b110;
      memory_array[1539] <= 3'b110;
      memory_array[1540] <= 3'b101;
      memory_array[1541] <= 3'b101;
      memory_array[1542] <= 3'b000;
      memory_array[1543] <= 3'b110;
      memory_array[1544] <= 3'b101;
      memory_array[1545] <= 3'b101;
      memory_array[1546] <= 3'b101;
      memory_array[1547] <= 3'b101;
      memory_array[1548] <= 3'b110;
      memory_array[1549] <= 3'b110;
      memory_array[1550] <= 3'b101;
      memory_array[1551] <= 3'b101;
      memory_array[1552] <= 3'b000;
      memory_array[1553] <= 3'b110;
      memory_array[1554] <= 3'b101;
      memory_array[1555] <= 3'b101;
      memory_array[1556] <= 3'b101;
      memory_array[1557] <= 3'b101;
      memory_array[1558] <= 3'b110;
      memory_array[1559] <= 3'b110;
      memory_array[1560] <= 3'b101;
      memory_array[1561] <= 3'b101;
      memory_array[1562] <= 3'b000;
      memory_array[1563] <= 3'b110;
      memory_array[1564] <= 3'b101;
      memory_array[1565] <= 3'b101;
      memory_array[1566] <= 3'b101;
      memory_array[1567] <= 3'b101;
      memory_array[1568] <= 3'b110;
      memory_array[1569] <= 3'b110;
      memory_array[1570] <= 3'b101;
      memory_array[1571] <= 3'b101;
      memory_array[1572] <= 3'b000;
      memory_array[1573] <= 3'b110;
      memory_array[1574] <= 3'b101;
      memory_array[1575] <= 3'b101;
      memory_array[1576] <= 3'b101;
      memory_array[1577] <= 3'b101;
      memory_array[1578] <= 3'b110;
      memory_array[1579] <= 3'b110;
      memory_array[1580] <= 3'b101;
      memory_array[1581] <= 3'b101;
      memory_array[1582] <= 3'b000;
      memory_array[1583] <= 3'b110;
      memory_array[1584] <= 3'b101;
      memory_array[1585] <= 3'b101;
      memory_array[1586] <= 3'b101;
      memory_array[1587] <= 3'b101;
      memory_array[1588] <= 3'b110;
      memory_array[1589] <= 3'b110;
      memory_array[1590] <= 3'b101;
      memory_array[1591] <= 3'b101;
      memory_array[1592] <= 3'b111;
      memory_array[1593] <= 3'b111;
      memory_array[1594] <= 3'b111;
      memory_array[1595] <= 3'b101;
      memory_array[1596] <= 3'b101;
      memory_array[1597] <= 3'b111;
      memory_array[1598] <= 3'b111;
      memory_array[1599] <= 3'b111;
      memory_array[1600] <= 3'b111;
      memory_array[1601] <= 3'b111;
      memory_array[1602] <= 3'b111;
      memory_array[1603] <= 3'b111;
      memory_array[1604] <= 3'b111;
      memory_array[1605] <= 3'b111;
      memory_array[1606] <= 3'b111;
      memory_array[1607] <= 3'b111;
      memory_array[1608] <= 3'b101;
      memory_array[1609] <= 3'b101;
      memory_array[1610] <= 3'b110;
      memory_array[1611] <= 3'b101;
      memory_array[1612] <= 3'b101;
      memory_array[1613] <= 3'b101;
      memory_array[1614] <= 3'b101;
      memory_array[1615] <= 3'b101;
      memory_array[1616] <= 3'b101;
      memory_array[1617] <= 3'b110;
      memory_array[1618] <= 3'b101;
      memory_array[1619] <= 3'b101;
      memory_array[1620] <= 3'b110;
      memory_array[1621] <= 3'b101;
      memory_array[1622] <= 3'b101;
      memory_array[1623] <= 3'b101;
      memory_array[1624] <= 3'b101;
      memory_array[1625] <= 3'b101;
      memory_array[1626] <= 3'b101;
      memory_array[1627] <= 3'b110;
      memory_array[1628] <= 3'b101;
      memory_array[1629] <= 3'b101;
      memory_array[1630] <= 3'b110;
      memory_array[1631] <= 3'b101;
      memory_array[1632] <= 3'b101;
      memory_array[1633] <= 3'b101;
      memory_array[1634] <= 3'b101;
      memory_array[1635] <= 3'b101;
      memory_array[1636] <= 3'b101;
      memory_array[1637] <= 3'b110;
      memory_array[1638] <= 3'b101;
      memory_array[1639] <= 3'b101;
      memory_array[1640] <= 3'b110;
      memory_array[1641] <= 3'b101;
      memory_array[1642] <= 3'b101;
      memory_array[1643] <= 3'b101;
      memory_array[1644] <= 3'b101;
      memory_array[1645] <= 3'b101;
      memory_array[1646] <= 3'b101;
      memory_array[1647] <= 3'b110;
      memory_array[1648] <= 3'b101;
      memory_array[1649] <= 3'b101;
      memory_array[1650] <= 3'b110;
      memory_array[1651] <= 3'b101;
      memory_array[1652] <= 3'b101;
      memory_array[1653] <= 3'b101;
      memory_array[1654] <= 3'b101;
      memory_array[1655] <= 3'b101;
      memory_array[1656] <= 3'b101;
      memory_array[1657] <= 3'b110;
      memory_array[1658] <= 3'b101;
      memory_array[1659] <= 3'b101;
      memory_array[1660] <= 3'b110;
      memory_array[1661] <= 3'b101;
      memory_array[1662] <= 3'b101;
      memory_array[1663] <= 3'b101;
      memory_array[1664] <= 3'b101;
      memory_array[1665] <= 3'b101;
      memory_array[1666] <= 3'b101;
      memory_array[1667] <= 3'b110;
      memory_array[1668] <= 3'b101;
      memory_array[1669] <= 3'b101;
      memory_array[1670] <= 3'b110;
      memory_array[1671] <= 3'b101;
      memory_array[1672] <= 3'b101;
      memory_array[1673] <= 3'b101;
      memory_array[1674] <= 3'b101;
      memory_array[1675] <= 3'b101;
      memory_array[1676] <= 3'b101;
      memory_array[1677] <= 3'b110;
      memory_array[1678] <= 3'b101;
      memory_array[1679] <= 3'b101;
      memory_array[1680] <= 3'b110;
      memory_array[1681] <= 3'b101;
      memory_array[1682] <= 3'b101;
      memory_array[1683] <= 3'b101;
      memory_array[1684] <= 3'b101;
      memory_array[1685] <= 3'b101;
      memory_array[1686] <= 3'b101;
      memory_array[1687] <= 3'b110;
      memory_array[1688] <= 3'b101;
      memory_array[1689] <= 3'b101;
      memory_array[1690] <= 3'b110;
      memory_array[1691] <= 3'b000;
      memory_array[1692] <= 3'b101;
      memory_array[1693] <= 3'b111;
      memory_array[1694] <= 3'b111;
      memory_array[1695] <= 3'b111;
      memory_array[1696] <= 3'b111;
      memory_array[1697] <= 3'b000;
      memory_array[1698] <= 3'b000;
      memory_array[1699] <= 3'b000;
      memory_array[1700] <= 3'b101;
      memory_array[1701] <= 3'b101;
      memory_array[1702] <= 3'b111;
      memory_array[1703] <= 3'b111;
      memory_array[1704] <= 3'b111;
      memory_array[1705] <= 3'b111;
      memory_array[1706] <= 3'b111;
      memory_array[1707] <= 3'b000;
      memory_array[1708] <= 3'b000;
      memory_array[1709] <= 3'b000;
      memory_array[1710] <= 3'b101;
      memory_array[1711] <= 3'b101;
      memory_array[1712] <= 3'b110;
      memory_array[1713] <= 3'b101;
      memory_array[1714] <= 3'b101;
      memory_array[1715] <= 3'b101;
      memory_array[1716] <= 3'b101;
      memory_array[1717] <= 3'b101;
      memory_array[1718] <= 3'b101;
      memory_array[1719] <= 3'b000;
      memory_array[1720] <= 3'b101;
      memory_array[1721] <= 3'b101;
      memory_array[1722] <= 3'b110;
      memory_array[1723] <= 3'b101;
      memory_array[1724] <= 3'b101;
      memory_array[1725] <= 3'b101;
      memory_array[1726] <= 3'b101;
      memory_array[1727] <= 3'b101;
      memory_array[1728] <= 3'b101;
      memory_array[1729] <= 3'b000;
      memory_array[1730] <= 3'b101;
      memory_array[1731] <= 3'b101;
      memory_array[1732] <= 3'b110;
      memory_array[1733] <= 3'b101;
      memory_array[1734] <= 3'b101;
      memory_array[1735] <= 3'b101;
      memory_array[1736] <= 3'b101;
      memory_array[1737] <= 3'b101;
      memory_array[1738] <= 3'b101;
      memory_array[1739] <= 3'b000;
      memory_array[1740] <= 3'b101;
      memory_array[1741] <= 3'b101;
      memory_array[1742] <= 3'b110;
      memory_array[1743] <= 3'b101;
      memory_array[1744] <= 3'b101;
      memory_array[1745] <= 3'b101;
      memory_array[1746] <= 3'b101;
      memory_array[1747] <= 3'b101;
      memory_array[1748] <= 3'b101;
      memory_array[1749] <= 3'b000;
      memory_array[1750] <= 3'b101;
      memory_array[1751] <= 3'b101;
      memory_array[1752] <= 3'b110;
      memory_array[1753] <= 3'b101;
      memory_array[1754] <= 3'b101;
      memory_array[1755] <= 3'b101;
      memory_array[1756] <= 3'b101;
      memory_array[1757] <= 3'b101;
      memory_array[1758] <= 3'b101;
      memory_array[1759] <= 3'b000;
      memory_array[1760] <= 3'b101;
      memory_array[1761] <= 3'b101;
      memory_array[1762] <= 3'b110;
      memory_array[1763] <= 3'b101;
      memory_array[1764] <= 3'b101;
      memory_array[1765] <= 3'b101;
      memory_array[1766] <= 3'b101;
      memory_array[1767] <= 3'b101;
      memory_array[1768] <= 3'b101;
      memory_array[1769] <= 3'b000;
      memory_array[1770] <= 3'b101;
      memory_array[1771] <= 3'b101;
      memory_array[1772] <= 3'b110;
      memory_array[1773] <= 3'b101;
      memory_array[1774] <= 3'b101;
      memory_array[1775] <= 3'b101;
      memory_array[1776] <= 3'b101;
      memory_array[1777] <= 3'b101;
      memory_array[1778] <= 3'b101;
      memory_array[1779] <= 3'b000;
      memory_array[1780] <= 3'b101;
      memory_array[1781] <= 3'b101;
      memory_array[1782] <= 3'b110;
      memory_array[1783] <= 3'b101;
      memory_array[1784] <= 3'b101;
      memory_array[1785] <= 3'b101;
      memory_array[1786] <= 3'b101;
      memory_array[1787] <= 3'b101;
      memory_array[1788] <= 3'b101;
      memory_array[1789] <= 3'b000;
      memory_array[1790] <= 3'b101;
      memory_array[1791] <= 3'b101;
      memory_array[1792] <= 3'b111;
      memory_array[1793] <= 3'b111;
      memory_array[1794] <= 3'b111;
      memory_array[1795] <= 3'b111;
      memory_array[1796] <= 3'b111;
      memory_array[1797] <= 3'b111;
      memory_array[1798] <= 3'b111;
      memory_array[1799] <= 3'b111;
      memory_array[1800] <= 3'b111;
      memory_array[1801] <= 3'b111;
      memory_array[1802] <= 3'b111;
      memory_array[1803] <= 3'b111;
      memory_array[1804] <= 3'b111;
      memory_array[1805] <= 3'b111;
      memory_array[1806] <= 3'b111;
      memory_array[1807] <= 3'b111;
      memory_array[1808] <= 3'b101;
      memory_array[1809] <= 3'b101;
      memory_array[1810] <= 3'b000;
      memory_array[1811] <= 3'b101;
      memory_array[1812] <= 3'b101;
      memory_array[1813] <= 3'b101;
      memory_array[1814] <= 3'b101;
      memory_array[1815] <= 3'b101;
      memory_array[1816] <= 3'b101;
      memory_array[1817] <= 3'b000;
      memory_array[1818] <= 3'b101;
      memory_array[1819] <= 3'b101;
      memory_array[1820] <= 3'b000;
      memory_array[1821] <= 3'b101;
      memory_array[1822] <= 3'b101;
      memory_array[1823] <= 3'b101;
      memory_array[1824] <= 3'b101;
      memory_array[1825] <= 3'b101;
      memory_array[1826] <= 3'b101;
      memory_array[1827] <= 3'b000;
      memory_array[1828] <= 3'b101;
      memory_array[1829] <= 3'b101;
      memory_array[1830] <= 3'b000;
      memory_array[1831] <= 3'b101;
      memory_array[1832] <= 3'b101;
      memory_array[1833] <= 3'b101;
      memory_array[1834] <= 3'b101;
      memory_array[1835] <= 3'b101;
      memory_array[1836] <= 3'b101;
      memory_array[1837] <= 3'b000;
      memory_array[1838] <= 3'b101;
      memory_array[1839] <= 3'b101;
      memory_array[1840] <= 3'b000;
      memory_array[1841] <= 3'b101;
      memory_array[1842] <= 3'b101;
      memory_array[1843] <= 3'b101;
      memory_array[1844] <= 3'b101;
      memory_array[1845] <= 3'b101;
      memory_array[1846] <= 3'b101;
      memory_array[1847] <= 3'b000;
      memory_array[1848] <= 3'b101;
      memory_array[1849] <= 3'b101;
      memory_array[1850] <= 3'b000;
      memory_array[1851] <= 3'b101;
      memory_array[1852] <= 3'b101;
      memory_array[1853] <= 3'b101;
      memory_array[1854] <= 3'b101;
      memory_array[1855] <= 3'b101;
      memory_array[1856] <= 3'b101;
      memory_array[1857] <= 3'b000;
      memory_array[1858] <= 3'b101;
      memory_array[1859] <= 3'b101;
      memory_array[1860] <= 3'b000;
      memory_array[1861] <= 3'b101;
      memory_array[1862] <= 3'b101;
      memory_array[1863] <= 3'b101;
      memory_array[1864] <= 3'b101;
      memory_array[1865] <= 3'b101;
      memory_array[1866] <= 3'b101;
      memory_array[1867] <= 3'b000;
      memory_array[1868] <= 3'b101;
      memory_array[1869] <= 3'b101;
      memory_array[1870] <= 3'b000;
      memory_array[1871] <= 3'b101;
      memory_array[1872] <= 3'b101;
      memory_array[1873] <= 3'b101;
      memory_array[1874] <= 3'b101;
      memory_array[1875] <= 3'b101;
      memory_array[1876] <= 3'b101;
      memory_array[1877] <= 3'b000;
      memory_array[1878] <= 3'b101;
      memory_array[1879] <= 3'b101;
      memory_array[1880] <= 3'b000;
      memory_array[1881] <= 3'b101;
      memory_array[1882] <= 3'b101;
      memory_array[1883] <= 3'b101;
      memory_array[1884] <= 3'b101;
      memory_array[1885] <= 3'b101;
      memory_array[1886] <= 3'b101;
      memory_array[1887] <= 3'b000;
      memory_array[1888] <= 3'b101;
      memory_array[1889] <= 3'b101;
      memory_array[1890] <= 3'b000;
      memory_array[1891] <= 3'b101;
      memory_array[1892] <= 3'b111;
      memory_array[1893] <= 3'b111;
      memory_array[1894] <= 3'b111;
      memory_array[1895] <= 3'b111;
      memory_array[1896] <= 3'b111;
      memory_array[1897] <= 3'b000;
      memory_array[1898] <= 3'b101;
      memory_array[1899] <= 3'b101;
      memory_array[1900] <= 3'b000;
      memory_array[1901] <= 3'b000;
      memory_array[1902] <= 3'b101;
      memory_array[1903] <= 3'b111;
      memory_array[1904] <= 3'b111;
      memory_array[1905] <= 3'b111;
      memory_array[1906] <= 3'b111;
      memory_array[1907] <= 3'b111;
      memory_array[1908] <= 3'b101;
      memory_array[1909] <= 3'b000;
      memory_array[1910] <= 3'b101;
      memory_array[1911] <= 3'b101;
      memory_array[1912] <= 3'b101;
      memory_array[1913] <= 3'b101;
      memory_array[1914] <= 3'b101;
      memory_array[1915] <= 3'b101;
      memory_array[1916] <= 3'b101;
      memory_array[1917] <= 3'b101;
      memory_array[1918] <= 3'b101;
      memory_array[1919] <= 3'b110;
      memory_array[1920] <= 3'b101;
      memory_array[1921] <= 3'b101;
      memory_array[1922] <= 3'b101;
      memory_array[1923] <= 3'b101;
      memory_array[1924] <= 3'b101;
      memory_array[1925] <= 3'b101;
      memory_array[1926] <= 3'b101;
      memory_array[1927] <= 3'b101;
      memory_array[1928] <= 3'b101;
      memory_array[1929] <= 3'b110;
      memory_array[1930] <= 3'b101;
      memory_array[1931] <= 3'b101;
      memory_array[1932] <= 3'b101;
      memory_array[1933] <= 3'b101;
      memory_array[1934] <= 3'b101;
      memory_array[1935] <= 3'b101;
      memory_array[1936] <= 3'b101;
      memory_array[1937] <= 3'b101;
      memory_array[1938] <= 3'b101;
      memory_array[1939] <= 3'b110;
      memory_array[1940] <= 3'b101;
      memory_array[1941] <= 3'b101;
      memory_array[1942] <= 3'b101;
      memory_array[1943] <= 3'b101;
      memory_array[1944] <= 3'b101;
      memory_array[1945] <= 3'b101;
      memory_array[1946] <= 3'b101;
      memory_array[1947] <= 3'b101;
      memory_array[1948] <= 3'b101;
      memory_array[1949] <= 3'b110;
      memory_array[1950] <= 3'b101;
      memory_array[1951] <= 3'b101;
      memory_array[1952] <= 3'b101;
      memory_array[1953] <= 3'b101;
      memory_array[1954] <= 3'b101;
      memory_array[1955] <= 3'b101;
      memory_array[1956] <= 3'b101;
      memory_array[1957] <= 3'b101;
      memory_array[1958] <= 3'b101;
      memory_array[1959] <= 3'b110;
      memory_array[1960] <= 3'b101;
      memory_array[1961] <= 3'b101;
      memory_array[1962] <= 3'b101;
      memory_array[1963] <= 3'b101;
      memory_array[1964] <= 3'b101;
      memory_array[1965] <= 3'b101;
      memory_array[1966] <= 3'b101;
      memory_array[1967] <= 3'b101;
      memory_array[1968] <= 3'b101;
      memory_array[1969] <= 3'b110;
      memory_array[1970] <= 3'b101;
      memory_array[1971] <= 3'b101;
      memory_array[1972] <= 3'b101;
      memory_array[1973] <= 3'b101;
      memory_array[1974] <= 3'b101;
      memory_array[1975] <= 3'b101;
      memory_array[1976] <= 3'b101;
      memory_array[1977] <= 3'b101;
      memory_array[1978] <= 3'b101;
      memory_array[1979] <= 3'b110;
      memory_array[1980] <= 3'b101;
      memory_array[1981] <= 3'b101;
      memory_array[1982] <= 3'b101;
      memory_array[1983] <= 3'b101;
      memory_array[1984] <= 3'b101;
      memory_array[1985] <= 3'b101;
      memory_array[1986] <= 3'b101;
      memory_array[1987] <= 3'b101;
      memory_array[1988] <= 3'b101;
      memory_array[1989] <= 3'b110;
      memory_array[1990] <= 3'b101;
      memory_array[1991] <= 3'b101;
      memory_array[1992] <= 3'b111;
      memory_array[1993] <= 3'b111;
      memory_array[1994] <= 3'b111;
      memory_array[1995] <= 3'b111;
      memory_array[1996] <= 3'b111;
      memory_array[1997] <= 3'b111;
      memory_array[1998] <= 3'b111;
      memory_array[1999] <= 3'b111;
      memory_array[2000] <= 3'b101;
      memory_array[2001] <= 3'b101;
      memory_array[2002] <= 3'b101;
      memory_array[2003] <= 3'b101;
      memory_array[2004] <= 3'b101;
      memory_array[2005] <= 3'b101;
      memory_array[2006] <= 3'b101;
      memory_array[2007] <= 3'b101;
      memory_array[2008] <= 3'b101;
      memory_array[2009] <= 3'b111;
      memory_array[2010] <= 3'b111;
      memory_array[2011] <= 3'b111;
      memory_array[2012] <= 3'b111;
      memory_array[2013] <= 3'b111;
      memory_array[2014] <= 3'b111;
      memory_array[2015] <= 3'b111;
      memory_array[2016] <= 3'b111;
      memory_array[2017] <= 3'b111;
      memory_array[2018] <= 3'b111;
      memory_array[2019] <= 3'b111;
      memory_array[2020] <= 3'b111;
      memory_array[2021] <= 3'b111;
      memory_array[2022] <= 3'b111;
      memory_array[2023] <= 3'b111;
      memory_array[2024] <= 3'b111;
      memory_array[2025] <= 3'b111;
      memory_array[2026] <= 3'b111;
      memory_array[2027] <= 3'b111;
      memory_array[2028] <= 3'b111;
      memory_array[2029] <= 3'b111;
      memory_array[2030] <= 3'b111;
      memory_array[2031] <= 3'b111;
      memory_array[2032] <= 3'b111;
      memory_array[2033] <= 3'b111;
      memory_array[2034] <= 3'b111;
      memory_array[2035] <= 3'b111;
      memory_array[2036] <= 3'b111;
      memory_array[2037] <= 3'b111;
      memory_array[2038] <= 3'b111;
      memory_array[2039] <= 3'b111;
      memory_array[2040] <= 3'b111;
      memory_array[2041] <= 3'b111;
      memory_array[2042] <= 3'b111;
      memory_array[2043] <= 3'b111;
      memory_array[2044] <= 3'b111;
      memory_array[2045] <= 3'b111;
      memory_array[2046] <= 3'b111;
      memory_array[2047] <= 3'b111;
      memory_array[2048] <= 3'b111;
      memory_array[2049] <= 3'b111;
      memory_array[2050] <= 3'b111;
      memory_array[2051] <= 3'b111;
      memory_array[2052] <= 3'b111;
      memory_array[2053] <= 3'b111;
      memory_array[2054] <= 3'b111;
      memory_array[2055] <= 3'b111;
      memory_array[2056] <= 3'b111;
      memory_array[2057] <= 3'b111;
      memory_array[2058] <= 3'b111;
      memory_array[2059] <= 3'b111;
      memory_array[2060] <= 3'b111;
      memory_array[2061] <= 3'b111;
      memory_array[2062] <= 3'b111;
      memory_array[2063] <= 3'b111;
      memory_array[2064] <= 3'b111;
      memory_array[2065] <= 3'b111;
      memory_array[2066] <= 3'b111;
      memory_array[2067] <= 3'b111;
      memory_array[2068] <= 3'b111;
      memory_array[2069] <= 3'b111;
      memory_array[2070] <= 3'b111;
      memory_array[2071] <= 3'b111;
      memory_array[2072] <= 3'b111;
      memory_array[2073] <= 3'b111;
      memory_array[2074] <= 3'b111;
      memory_array[2075] <= 3'b111;
      memory_array[2076] <= 3'b111;
      memory_array[2077] <= 3'b111;
      memory_array[2078] <= 3'b111;
      memory_array[2079] <= 3'b111;
      memory_array[2080] <= 3'b111;
      memory_array[2081] <= 3'b111;
      memory_array[2082] <= 3'b111;
      memory_array[2083] <= 3'b111;
      memory_array[2084] <= 3'b111;
      memory_array[2085] <= 3'b111;
      memory_array[2086] <= 3'b101;
      memory_array[2087] <= 3'b000;
      memory_array[2088] <= 3'b000;
      memory_array[2089] <= 3'b000;
      memory_array[2090] <= 3'b101;
      memory_array[2091] <= 3'b111;
      memory_array[2092] <= 3'b111;
      memory_array[2093] <= 3'b111;
      memory_array[2094] <= 3'b111;
      memory_array[2095] <= 3'b111;
      memory_array[2096] <= 3'b101;
      memory_array[2097] <= 3'b101;
      memory_array[2098] <= 3'b000;
      memory_array[2099] <= 3'b000;
      memory_array[2100] <= 3'b101;
      memory_array[2101] <= 3'b101;
      memory_array[2102] <= 3'b000;
      memory_array[2103] <= 3'b101;
      memory_array[2104] <= 3'b111;
      memory_array[2105] <= 3'b111;
      memory_array[2106] <= 3'b111;
      memory_array[2107] <= 3'b111;
      memory_array[2108] <= 3'b111;
      memory_array[2109] <= 3'b101;
      memory_array[2110] <= 3'b000;
      memory_array[2111] <= 3'b000;
      memory_array[2112] <= 3'b101;
      memory_array[2113] <= 3'b101;
      memory_array[2114] <= 3'b111;
      memory_array[2115] <= 3'b111;
      memory_array[2116] <= 3'b111;
      memory_array[2117] <= 3'b111;
      memory_array[2118] <= 3'b111;
      memory_array[2119] <= 3'b111;
      memory_array[2120] <= 3'b111;
      memory_array[2121] <= 3'b111;
      memory_array[2122] <= 3'b111;
      memory_array[2123] <= 3'b111;
      memory_array[2124] <= 3'b111;
      memory_array[2125] <= 3'b111;
      memory_array[2126] <= 3'b111;
      memory_array[2127] <= 3'b111;
      memory_array[2128] <= 3'b111;
      memory_array[2129] <= 3'b111;
      memory_array[2130] <= 3'b111;
      memory_array[2131] <= 3'b111;
      memory_array[2132] <= 3'b111;
      memory_array[2133] <= 3'b111;
      memory_array[2134] <= 3'b111;
      memory_array[2135] <= 3'b111;
      memory_array[2136] <= 3'b111;
      memory_array[2137] <= 3'b111;
      memory_array[2138] <= 3'b111;
      memory_array[2139] <= 3'b111;
      memory_array[2140] <= 3'b111;
      memory_array[2141] <= 3'b111;
      memory_array[2142] <= 3'b111;
      memory_array[2143] <= 3'b111;
      memory_array[2144] <= 3'b111;
      memory_array[2145] <= 3'b111;
      memory_array[2146] <= 3'b111;
      memory_array[2147] <= 3'b111;
      memory_array[2148] <= 3'b111;
      memory_array[2149] <= 3'b111;
      memory_array[2150] <= 3'b111;
      memory_array[2151] <= 3'b111;
      memory_array[2152] <= 3'b111;
      memory_array[2153] <= 3'b111;
      memory_array[2154] <= 3'b111;
      memory_array[2155] <= 3'b111;
      memory_array[2156] <= 3'b111;
      memory_array[2157] <= 3'b111;
      memory_array[2158] <= 3'b111;
      memory_array[2159] <= 3'b111;
      memory_array[2160] <= 3'b111;
      memory_array[2161] <= 3'b111;
      memory_array[2162] <= 3'b111;
      memory_array[2163] <= 3'b111;
      memory_array[2164] <= 3'b111;
      memory_array[2165] <= 3'b111;
      memory_array[2166] <= 3'b111;
      memory_array[2167] <= 3'b111;
      memory_array[2168] <= 3'b111;
      memory_array[2169] <= 3'b111;
      memory_array[2170] <= 3'b111;
      memory_array[2171] <= 3'b111;
      memory_array[2172] <= 3'b111;
      memory_array[2173] <= 3'b111;
      memory_array[2174] <= 3'b111;
      memory_array[2175] <= 3'b111;
      memory_array[2176] <= 3'b111;
      memory_array[2177] <= 3'b111;
      memory_array[2178] <= 3'b111;
      memory_array[2179] <= 3'b111;
      memory_array[2180] <= 3'b111;
      memory_array[2181] <= 3'b111;
      memory_array[2182] <= 3'b111;
      memory_array[2183] <= 3'b111;
      memory_array[2184] <= 3'b111;
      memory_array[2185] <= 3'b111;
      memory_array[2186] <= 3'b111;
      memory_array[2187] <= 3'b111;
      memory_array[2188] <= 3'b111;
      memory_array[2189] <= 3'b111;
      memory_array[2190] <= 3'b111;
      memory_array[2191] <= 3'b101;
      memory_array[2192] <= 3'b101;
      memory_array[2193] <= 3'b101;
      memory_array[2194] <= 3'b101;
      memory_array[2195] <= 3'b101;
      memory_array[2196] <= 3'b101;
      memory_array[2197] <= 3'b101;
      memory_array[2198] <= 3'b101;
      memory_array[2199] <= 3'b101;
      memory_array[2200] <= 3'b101;
      memory_array[2201] <= 3'b101;
      memory_array[2202] <= 3'b101;
      memory_array[2203] <= 3'b101;
      memory_array[2204] <= 3'b101;
      memory_array[2205] <= 3'b101;
      memory_array[2206] <= 3'b101;
      memory_array[2207] <= 3'b101;
      memory_array[2208] <= 3'b101;
      memory_array[2209] <= 3'b000;
      memory_array[2210] <= 3'b000;
      memory_array[2211] <= 3'b000;
      memory_array[2212] <= 3'b000;
      memory_array[2213] <= 3'b000;
      memory_array[2214] <= 3'b000;
      memory_array[2215] <= 3'b000;
      memory_array[2216] <= 3'b000;
      memory_array[2217] <= 3'b000;
      memory_array[2218] <= 3'b000;
      memory_array[2219] <= 3'b000;
      memory_array[2220] <= 3'b000;
      memory_array[2221] <= 3'b000;
      memory_array[2222] <= 3'b000;
      memory_array[2223] <= 3'b000;
      memory_array[2224] <= 3'b000;
      memory_array[2225] <= 3'b000;
      memory_array[2226] <= 3'b000;
      memory_array[2227] <= 3'b000;
      memory_array[2228] <= 3'b000;
      memory_array[2229] <= 3'b000;
      memory_array[2230] <= 3'b000;
      memory_array[2231] <= 3'b000;
      memory_array[2232] <= 3'b000;
      memory_array[2233] <= 3'b000;
      memory_array[2234] <= 3'b000;
      memory_array[2235] <= 3'b000;
      memory_array[2236] <= 3'b000;
      memory_array[2237] <= 3'b000;
      memory_array[2238] <= 3'b000;
      memory_array[2239] <= 3'b000;
      memory_array[2240] <= 3'b000;
      memory_array[2241] <= 3'b000;
      memory_array[2242] <= 3'b000;
      memory_array[2243] <= 3'b000;
      memory_array[2244] <= 3'b000;
      memory_array[2245] <= 3'b000;
      memory_array[2246] <= 3'b000;
      memory_array[2247] <= 3'b000;
      memory_array[2248] <= 3'b000;
      memory_array[2249] <= 3'b000;
      memory_array[2250] <= 3'b000;
      memory_array[2251] <= 3'b000;
      memory_array[2252] <= 3'b000;
      memory_array[2253] <= 3'b000;
      memory_array[2254] <= 3'b000;
      memory_array[2255] <= 3'b000;
      memory_array[2256] <= 3'b000;
      memory_array[2257] <= 3'b000;
      memory_array[2258] <= 3'b000;
      memory_array[2259] <= 3'b000;
      memory_array[2260] <= 3'b000;
      memory_array[2261] <= 3'b000;
      memory_array[2262] <= 3'b000;
      memory_array[2263] <= 3'b000;
      memory_array[2264] <= 3'b000;
      memory_array[2265] <= 3'b000;
      memory_array[2266] <= 3'b000;
      memory_array[2267] <= 3'b000;
      memory_array[2268] <= 3'b000;
      memory_array[2269] <= 3'b000;
      memory_array[2270] <= 3'b000;
      memory_array[2271] <= 3'b000;
      memory_array[2272] <= 3'b000;
      memory_array[2273] <= 3'b000;
      memory_array[2274] <= 3'b000;
      memory_array[2275] <= 3'b000;
      memory_array[2276] <= 3'b000;
      memory_array[2277] <= 3'b000;
      memory_array[2278] <= 3'b000;
      memory_array[2279] <= 3'b000;
      memory_array[2280] <= 3'b000;
      memory_array[2281] <= 3'b000;
      memory_array[2282] <= 3'b000;
      memory_array[2283] <= 3'b000;
      memory_array[2284] <= 3'b000;
      memory_array[2285] <= 3'b000;
      memory_array[2286] <= 3'b101;
      memory_array[2287] <= 3'b111;
      memory_array[2288] <= 3'b111;
      memory_array[2289] <= 3'b111;
      memory_array[2290] <= 3'b111;
      memory_array[2291] <= 3'b111;
      memory_array[2292] <= 3'b111;
      memory_array[2293] <= 3'b111;
      memory_array[2294] <= 3'b111;
      memory_array[2295] <= 3'b101;
      memory_array[2296] <= 3'b101;
      memory_array[2297] <= 3'b101;
      memory_array[2298] <= 3'b000;
      memory_array[2299] <= 3'b000;
      memory_array[2300] <= 3'b101;
      memory_array[2301] <= 3'b101;
      memory_array[2302] <= 3'b101;
      memory_array[2303] <= 3'b000;
      memory_array[2304] <= 3'b101;
      memory_array[2305] <= 3'b111;
      memory_array[2306] <= 3'b111;
      memory_array[2307] <= 3'b111;
      memory_array[2308] <= 3'b111;
      memory_array[2309] <= 3'b111;
      memory_array[2310] <= 3'b111;
      memory_array[2311] <= 3'b111;
      memory_array[2312] <= 3'b111;
      memory_array[2313] <= 3'b101;
      memory_array[2314] <= 3'b000;
      memory_array[2315] <= 3'b000;
      memory_array[2316] <= 3'b000;
      memory_array[2317] <= 3'b000;
      memory_array[2318] <= 3'b000;
      memory_array[2319] <= 3'b000;
      memory_array[2320] <= 3'b000;
      memory_array[2321] <= 3'b000;
      memory_array[2322] <= 3'b000;
      memory_array[2323] <= 3'b000;
      memory_array[2324] <= 3'b000;
      memory_array[2325] <= 3'b000;
      memory_array[2326] <= 3'b000;
      memory_array[2327] <= 3'b000;
      memory_array[2328] <= 3'b000;
      memory_array[2329] <= 3'b000;
      memory_array[2330] <= 3'b000;
      memory_array[2331] <= 3'b000;
      memory_array[2332] <= 3'b000;
      memory_array[2333] <= 3'b000;
      memory_array[2334] <= 3'b000;
      memory_array[2335] <= 3'b000;
      memory_array[2336] <= 3'b000;
      memory_array[2337] <= 3'b000;
      memory_array[2338] <= 3'b000;
      memory_array[2339] <= 3'b000;
      memory_array[2340] <= 3'b000;
      memory_array[2341] <= 3'b000;
      memory_array[2342] <= 3'b000;
      memory_array[2343] <= 3'b000;
      memory_array[2344] <= 3'b000;
      memory_array[2345] <= 3'b000;
      memory_array[2346] <= 3'b000;
      memory_array[2347] <= 3'b000;
      memory_array[2348] <= 3'b000;
      memory_array[2349] <= 3'b000;
      memory_array[2350] <= 3'b000;
      memory_array[2351] <= 3'b000;
      memory_array[2352] <= 3'b000;
      memory_array[2353] <= 3'b000;
      memory_array[2354] <= 3'b000;
      memory_array[2355] <= 3'b000;
      memory_array[2356] <= 3'b000;
      memory_array[2357] <= 3'b000;
      memory_array[2358] <= 3'b000;
      memory_array[2359] <= 3'b000;
      memory_array[2360] <= 3'b000;
      memory_array[2361] <= 3'b000;
      memory_array[2362] <= 3'b000;
      memory_array[2363] <= 3'b000;
      memory_array[2364] <= 3'b000;
      memory_array[2365] <= 3'b000;
      memory_array[2366] <= 3'b000;
      memory_array[2367] <= 3'b000;
      memory_array[2368] <= 3'b000;
      memory_array[2369] <= 3'b000;
      memory_array[2370] <= 3'b000;
      memory_array[2371] <= 3'b000;
      memory_array[2372] <= 3'b000;
      memory_array[2373] <= 3'b000;
      memory_array[2374] <= 3'b000;
      memory_array[2375] <= 3'b000;
      memory_array[2376] <= 3'b000;
      memory_array[2377] <= 3'b000;
      memory_array[2378] <= 3'b000;
      memory_array[2379] <= 3'b000;
      memory_array[2380] <= 3'b000;
      memory_array[2381] <= 3'b000;
      memory_array[2382] <= 3'b000;
      memory_array[2383] <= 3'b000;
      memory_array[2384] <= 3'b000;
      memory_array[2385] <= 3'b000;
      memory_array[2386] <= 3'b000;
      memory_array[2387] <= 3'b000;
      memory_array[2388] <= 3'b000;
      memory_array[2389] <= 3'b000;
      memory_array[2390] <= 3'b000;
      memory_array[2391] <= 3'b101;
      memory_array[2392] <= 3'b101;
      memory_array[2393] <= 3'b101;
      memory_array[2394] <= 3'b101;
      memory_array[2395] <= 3'b101;
      memory_array[2396] <= 3'b101;
      memory_array[2397] <= 3'b101;
      memory_array[2398] <= 3'b101;
      memory_array[2399] <= 3'b101;
      memory_array[2400] <= 3'b000;
      memory_array[2401] <= 3'b000;
      memory_array[2402] <= 3'b000;
      memory_array[2403] <= 3'b110;
      memory_array[2404] <= 3'b110;
      memory_array[2405] <= 3'b000;
      memory_array[2406] <= 3'b000;
      memory_array[2407] <= 3'b000;
      memory_array[2408] <= 3'b101;
      memory_array[2409] <= 3'b000;
      memory_array[2410] <= 3'b000;
      memory_array[2411] <= 3'b000;
      memory_array[2412] <= 3'b000;
      memory_array[2413] <= 3'b000;
      memory_array[2414] <= 3'b000;
      memory_array[2415] <= 3'b000;
      memory_array[2416] <= 3'b000;
      memory_array[2417] <= 3'b000;
      memory_array[2418] <= 3'b000;
      memory_array[2419] <= 3'b000;
      memory_array[2420] <= 3'b000;
      memory_array[2421] <= 3'b000;
      memory_array[2422] <= 3'b000;
      memory_array[2423] <= 3'b000;
      memory_array[2424] <= 3'b000;
      memory_array[2425] <= 3'b000;
      memory_array[2426] <= 3'b000;
      memory_array[2427] <= 3'b000;
      memory_array[2428] <= 3'b000;
      memory_array[2429] <= 3'b000;
      memory_array[2430] <= 3'b000;
      memory_array[2431] <= 3'b000;
      memory_array[2432] <= 3'b000;
      memory_array[2433] <= 3'b000;
      memory_array[2434] <= 3'b000;
      memory_array[2435] <= 3'b000;
      memory_array[2436] <= 3'b000;
      memory_array[2437] <= 3'b000;
      memory_array[2438] <= 3'b000;
      memory_array[2439] <= 3'b000;
      memory_array[2440] <= 3'b000;
      memory_array[2441] <= 3'b000;
      memory_array[2442] <= 3'b000;
      memory_array[2443] <= 3'b000;
      memory_array[2444] <= 3'b000;
      memory_array[2445] <= 3'b000;
      memory_array[2446] <= 3'b000;
      memory_array[2447] <= 3'b000;
      memory_array[2448] <= 3'b000;
      memory_array[2449] <= 3'b000;
      memory_array[2450] <= 3'b000;
      memory_array[2451] <= 3'b000;
      memory_array[2452] <= 3'b000;
      memory_array[2453] <= 3'b000;
      memory_array[2454] <= 3'b000;
      memory_array[2455] <= 3'b000;
      memory_array[2456] <= 3'b000;
      memory_array[2457] <= 3'b000;
      memory_array[2458] <= 3'b000;
      memory_array[2459] <= 3'b000;
      memory_array[2460] <= 3'b000;
      memory_array[2461] <= 3'b000;
      memory_array[2462] <= 3'b000;
      memory_array[2463] <= 3'b000;
      memory_array[2464] <= 3'b000;
      memory_array[2465] <= 3'b000;
      memory_array[2466] <= 3'b000;
      memory_array[2467] <= 3'b000;
      memory_array[2468] <= 3'b000;
      memory_array[2469] <= 3'b000;
      memory_array[2470] <= 3'b000;
      memory_array[2471] <= 3'b000;
      memory_array[2472] <= 3'b000;
      memory_array[2473] <= 3'b000;
      memory_array[2474] <= 3'b000;
      memory_array[2475] <= 3'b000;
      memory_array[2476] <= 3'b000;
      memory_array[2477] <= 3'b000;
      memory_array[2478] <= 3'b000;
      memory_array[2479] <= 3'b000;
      memory_array[2480] <= 3'b000;
      memory_array[2481] <= 3'b000;
      memory_array[2482] <= 3'b101;
      memory_array[2483] <= 3'b101;
      memory_array[2484] <= 3'b111;
      memory_array[2485] <= 3'b111;
      memory_array[2486] <= 3'b111;
      memory_array[2487] <= 3'b111;
      memory_array[2488] <= 3'b111;
      memory_array[2489] <= 3'b111;
      memory_array[2490] <= 3'b111;
      memory_array[2491] <= 3'b111;
      memory_array[2492] <= 3'b111;
      memory_array[2493] <= 3'b111;
      memory_array[2494] <= 3'b000;
      memory_array[2495] <= 3'b000;
      memory_array[2496] <= 3'b000;
      memory_array[2497] <= 3'b000;
      memory_array[2498] <= 3'b101;
      memory_array[2499] <= 3'b101;
      memory_array[2500] <= 3'b000;
      memory_array[2501] <= 3'b000;
      memory_array[2502] <= 3'b000;
      memory_array[2503] <= 3'b101;
      memory_array[2504] <= 3'b000;
      memory_array[2505] <= 3'b000;
      memory_array[2506] <= 3'b111;
      memory_array[2507] <= 3'b111;
      memory_array[2508] <= 3'b111;
      memory_array[2509] <= 3'b111;
      memory_array[2510] <= 3'b111;
      memory_array[2511] <= 3'b111;
      memory_array[2512] <= 3'b111;
      memory_array[2513] <= 3'b111;
      memory_array[2514] <= 3'b111;
      memory_array[2515] <= 3'b111;
      memory_array[2516] <= 3'b101;
      memory_array[2517] <= 3'b000;
      memory_array[2518] <= 3'b000;
      memory_array[2519] <= 3'b000;
      memory_array[2520] <= 3'b000;
      memory_array[2521] <= 3'b000;
      memory_array[2522] <= 3'b000;
      memory_array[2523] <= 3'b000;
      memory_array[2524] <= 3'b000;
      memory_array[2525] <= 3'b000;
      memory_array[2526] <= 3'b000;
      memory_array[2527] <= 3'b000;
      memory_array[2528] <= 3'b000;
      memory_array[2529] <= 3'b000;
      memory_array[2530] <= 3'b000;
      memory_array[2531] <= 3'b000;
      memory_array[2532] <= 3'b000;
      memory_array[2533] <= 3'b000;
      memory_array[2534] <= 3'b000;
      memory_array[2535] <= 3'b000;
      memory_array[2536] <= 3'b000;
      memory_array[2537] <= 3'b000;
      memory_array[2538] <= 3'b000;
      memory_array[2539] <= 3'b000;
      memory_array[2540] <= 3'b000;
      memory_array[2541] <= 3'b000;
      memory_array[2542] <= 3'b000;
      memory_array[2543] <= 3'b000;
      memory_array[2544] <= 3'b000;
      memory_array[2545] <= 3'b000;
      memory_array[2546] <= 3'b000;
      memory_array[2547] <= 3'b000;
      memory_array[2548] <= 3'b000;
      memory_array[2549] <= 3'b000;
      memory_array[2550] <= 3'b000;
      memory_array[2551] <= 3'b000;
      memory_array[2552] <= 3'b000;
      memory_array[2553] <= 3'b000;
      memory_array[2554] <= 3'b000;
      memory_array[2555] <= 3'b000;
      memory_array[2556] <= 3'b000;
      memory_array[2557] <= 3'b000;
      memory_array[2558] <= 3'b000;
      memory_array[2559] <= 3'b000;
      memory_array[2560] <= 3'b000;
      memory_array[2561] <= 3'b000;
      memory_array[2562] <= 3'b000;
      memory_array[2563] <= 3'b000;
      memory_array[2564] <= 3'b000;
      memory_array[2565] <= 3'b000;
      memory_array[2566] <= 3'b000;
      memory_array[2567] <= 3'b000;
      memory_array[2568] <= 3'b000;
      memory_array[2569] <= 3'b000;
      memory_array[2570] <= 3'b000;
      memory_array[2571] <= 3'b000;
      memory_array[2572] <= 3'b000;
      memory_array[2573] <= 3'b000;
      memory_array[2574] <= 3'b000;
      memory_array[2575] <= 3'b000;
      memory_array[2576] <= 3'b000;
      memory_array[2577] <= 3'b000;
      memory_array[2578] <= 3'b000;
      memory_array[2579] <= 3'b000;
      memory_array[2580] <= 3'b000;
      memory_array[2581] <= 3'b000;
      memory_array[2582] <= 3'b000;
      memory_array[2583] <= 3'b000;
      memory_array[2584] <= 3'b000;
      memory_array[2585] <= 3'b000;
      memory_array[2586] <= 3'b000;
      memory_array[2587] <= 3'b000;
      memory_array[2588] <= 3'b000;
      memory_array[2589] <= 3'b000;
      memory_array[2590] <= 3'b000;
      memory_array[2591] <= 3'b101;
      memory_array[2592] <= 3'b000;
      memory_array[2593] <= 3'b110;
      memory_array[2594] <= 3'b110;
      memory_array[2595] <= 3'b000;
      memory_array[2596] <= 3'b000;
      memory_array[2597] <= 3'b000;
      memory_array[2598] <= 3'b110;
      memory_array[2599] <= 3'b110;
      memory_array[2600] <= 3'b101;
      memory_array[2601] <= 3'b110;
      memory_array[2602] <= 3'b110;
      memory_array[2603] <= 3'b000;
      memory_array[2604] <= 3'b000;
      memory_array[2605] <= 3'b110;
      memory_array[2606] <= 3'b110;
      memory_array[2607] <= 3'b101;
      memory_array[2608] <= 3'b101;
      memory_array[2609] <= 3'b000;
      memory_array[2610] <= 3'b000;
      memory_array[2611] <= 3'b000;
      memory_array[2612] <= 3'b000;
      memory_array[2613] <= 3'b000;
      memory_array[2614] <= 3'b000;
      memory_array[2615] <= 3'b000;
      memory_array[2616] <= 3'b000;
      memory_array[2617] <= 3'b000;
      memory_array[2618] <= 3'b000;
      memory_array[2619] <= 3'b000;
      memory_array[2620] <= 3'b000;
      memory_array[2621] <= 3'b000;
      memory_array[2622] <= 3'b000;
      memory_array[2623] <= 3'b000;
      memory_array[2624] <= 3'b000;
      memory_array[2625] <= 3'b000;
      memory_array[2626] <= 3'b000;
      memory_array[2627] <= 3'b000;
      memory_array[2628] <= 3'b000;
      memory_array[2629] <= 3'b000;
      memory_array[2630] <= 3'b000;
      memory_array[2631] <= 3'b000;
      memory_array[2632] <= 3'b000;
      memory_array[2633] <= 3'b000;
      memory_array[2634] <= 3'b000;
      memory_array[2635] <= 3'b000;
      memory_array[2636] <= 3'b000;
      memory_array[2637] <= 3'b000;
      memory_array[2638] <= 3'b000;
      memory_array[2639] <= 3'b000;
      memory_array[2640] <= 3'b000;
      memory_array[2641] <= 3'b000;
      memory_array[2642] <= 3'b000;
      memory_array[2643] <= 3'b000;
      memory_array[2644] <= 3'b000;
      memory_array[2645] <= 3'b000;
      memory_array[2646] <= 3'b000;
      memory_array[2647] <= 3'b000;
      memory_array[2648] <= 3'b000;
      memory_array[2649] <= 3'b000;
      memory_array[2650] <= 3'b000;
      memory_array[2651] <= 3'b000;
      memory_array[2652] <= 3'b000;
      memory_array[2653] <= 3'b000;
      memory_array[2654] <= 3'b000;
      memory_array[2655] <= 3'b000;
      memory_array[2656] <= 3'b000;
      memory_array[2657] <= 3'b000;
      memory_array[2658] <= 3'b000;
      memory_array[2659] <= 3'b000;
      memory_array[2660] <= 3'b000;
      memory_array[2661] <= 3'b000;
      memory_array[2662] <= 3'b000;
      memory_array[2663] <= 3'b000;
      memory_array[2664] <= 3'b000;
      memory_array[2665] <= 3'b000;
      memory_array[2666] <= 3'b000;
      memory_array[2667] <= 3'b000;
      memory_array[2668] <= 3'b000;
      memory_array[2669] <= 3'b000;
      memory_array[2670] <= 3'b000;
      memory_array[2671] <= 3'b000;
      memory_array[2672] <= 3'b000;
      memory_array[2673] <= 3'b000;
      memory_array[2674] <= 3'b000;
      memory_array[2675] <= 3'b000;
      memory_array[2676] <= 3'b000;
      memory_array[2677] <= 3'b000;
      memory_array[2678] <= 3'b000;
      memory_array[2679] <= 3'b000;
      memory_array[2680] <= 3'b000;
      memory_array[2681] <= 3'b111;
      memory_array[2682] <= 3'b111;
      memory_array[2683] <= 3'b111;
      memory_array[2684] <= 3'b111;
      memory_array[2685] <= 3'b111;
      memory_array[2686] <= 3'b111;
      memory_array[2687] <= 3'b111;
      memory_array[2688] <= 3'b111;
      memory_array[2689] <= 3'b111;
      memory_array[2690] <= 3'b111;
      memory_array[2691] <= 3'b111;
      memory_array[2692] <= 3'b101;
      memory_array[2693] <= 3'b000;
      memory_array[2694] <= 3'b000;
      memory_array[2695] <= 3'b101;
      memory_array[2696] <= 3'b101;
      memory_array[2697] <= 3'b101;
      memory_array[2698] <= 3'b000;
      memory_array[2699] <= 3'b000;
      memory_array[2700] <= 3'b101;
      memory_array[2701] <= 3'b101;
      memory_array[2702] <= 3'b101;
      memory_array[2703] <= 3'b000;
      memory_array[2704] <= 3'b000;
      memory_array[2705] <= 3'b101;
      memory_array[2706] <= 3'b000;
      memory_array[2707] <= 3'b111;
      memory_array[2708] <= 3'b111;
      memory_array[2709] <= 3'b111;
      memory_array[2710] <= 3'b111;
      memory_array[2711] <= 3'b111;
      memory_array[2712] <= 3'b111;
      memory_array[2713] <= 3'b111;
      memory_array[2714] <= 3'b111;
      memory_array[2715] <= 3'b111;
      memory_array[2716] <= 3'b111;
      memory_array[2717] <= 3'b111;
      memory_array[2718] <= 3'b111;
      memory_array[2719] <= 3'b000;
      memory_array[2720] <= 3'b000;
      memory_array[2721] <= 3'b000;
      memory_array[2722] <= 3'b000;
      memory_array[2723] <= 3'b000;
      memory_array[2724] <= 3'b000;
      memory_array[2725] <= 3'b000;
      memory_array[2726] <= 3'b000;
      memory_array[2727] <= 3'b000;
      memory_array[2728] <= 3'b000;
      memory_array[2729] <= 3'b000;
      memory_array[2730] <= 3'b000;
      memory_array[2731] <= 3'b000;
      memory_array[2732] <= 3'b000;
      memory_array[2733] <= 3'b000;
      memory_array[2734] <= 3'b000;
      memory_array[2735] <= 3'b000;
      memory_array[2736] <= 3'b000;
      memory_array[2737] <= 3'b000;
      memory_array[2738] <= 3'b000;
      memory_array[2739] <= 3'b000;
      memory_array[2740] <= 3'b000;
      memory_array[2741] <= 3'b000;
      memory_array[2742] <= 3'b000;
      memory_array[2743] <= 3'b000;
      memory_array[2744] <= 3'b000;
      memory_array[2745] <= 3'b000;
      memory_array[2746] <= 3'b000;
      memory_array[2747] <= 3'b000;
      memory_array[2748] <= 3'b000;
      memory_array[2749] <= 3'b000;
      memory_array[2750] <= 3'b000;
      memory_array[2751] <= 3'b000;
      memory_array[2752] <= 3'b000;
      memory_array[2753] <= 3'b000;
      memory_array[2754] <= 3'b000;
      memory_array[2755] <= 3'b000;
      memory_array[2756] <= 3'b000;
      memory_array[2757] <= 3'b000;
      memory_array[2758] <= 3'b000;
      memory_array[2759] <= 3'b000;
      memory_array[2760] <= 3'b000;
      memory_array[2761] <= 3'b000;
      memory_array[2762] <= 3'b000;
      memory_array[2763] <= 3'b000;
      memory_array[2764] <= 3'b000;
      memory_array[2765] <= 3'b000;
      memory_array[2766] <= 3'b000;
      memory_array[2767] <= 3'b000;
      memory_array[2768] <= 3'b000;
      memory_array[2769] <= 3'b000;
      memory_array[2770] <= 3'b000;
      memory_array[2771] <= 3'b000;
      memory_array[2772] <= 3'b000;
      memory_array[2773] <= 3'b000;
      memory_array[2774] <= 3'b000;
      memory_array[2775] <= 3'b000;
      memory_array[2776] <= 3'b000;
      memory_array[2777] <= 3'b000;
      memory_array[2778] <= 3'b000;
      memory_array[2779] <= 3'b000;
      memory_array[2780] <= 3'b000;
      memory_array[2781] <= 3'b000;
      memory_array[2782] <= 3'b000;
      memory_array[2783] <= 3'b000;
      memory_array[2784] <= 3'b000;
      memory_array[2785] <= 3'b000;
      memory_array[2786] <= 3'b000;
      memory_array[2787] <= 3'b000;
      memory_array[2788] <= 3'b000;
      memory_array[2789] <= 3'b000;
      memory_array[2790] <= 3'b000;
      memory_array[2791] <= 3'b101;
      memory_array[2792] <= 3'b110;
      memory_array[2793] <= 3'b000;
      memory_array[2794] <= 3'b000;
      memory_array[2795] <= 3'b110;
      memory_array[2796] <= 3'b110;
      memory_array[2797] <= 3'b110;
      memory_array[2798] <= 3'b000;
      memory_array[2799] <= 3'b101;
      memory_array[2800] <= 3'b101;
      memory_array[2801] <= 3'b101;
      memory_array[2802] <= 3'b110;
      memory_array[2803] <= 3'b101;
      memory_array[2804] <= 3'b101;
      memory_array[2805] <= 3'b110;
      memory_array[2806] <= 3'b101;
      memory_array[2807] <= 3'b101;
      memory_array[2808] <= 3'b101;
      memory_array[2809] <= 3'b000;
      memory_array[2810] <= 3'b000;
      memory_array[2811] <= 3'b101;
      memory_array[2812] <= 3'b000;
      memory_array[2813] <= 3'b101;
      memory_array[2814] <= 3'b101;
      memory_array[2815] <= 3'b000;
      memory_array[2816] <= 3'b101;
      memory_array[2817] <= 3'b110;
      memory_array[2818] <= 3'b000;
      memory_array[2819] <= 3'b000;
      memory_array[2820] <= 3'b110;
      memory_array[2821] <= 3'b000;
      memory_array[2822] <= 3'b000;
      memory_array[2823] <= 3'b000;
      memory_array[2824] <= 3'b000;
      memory_array[2825] <= 3'b110;
      memory_array[2826] <= 3'b000;
      memory_array[2827] <= 3'b101;
      memory_array[2828] <= 3'b000;
      memory_array[2829] <= 3'b000;
      memory_array[2830] <= 3'b110;
      memory_array[2831] <= 3'b110;
      memory_array[2832] <= 3'b110;
      memory_array[2833] <= 3'b000;
      memory_array[2834] <= 3'b000;
      memory_array[2835] <= 3'b110;
      memory_array[2836] <= 3'b000;
      memory_array[2837] <= 3'b000;
      memory_array[2838] <= 3'b000;
      memory_array[2839] <= 3'b000;
      memory_array[2840] <= 3'b101;
      memory_array[2841] <= 3'b000;
      memory_array[2842] <= 3'b110;
      memory_array[2843] <= 3'b000;
      memory_array[2844] <= 3'b000;
      memory_array[2845] <= 3'b110;
      memory_array[2846] <= 3'b101;
      memory_array[2847] <= 3'b000;
      memory_array[2848] <= 3'b101;
      memory_array[2849] <= 3'b101;
      memory_array[2850] <= 3'b000;
      memory_array[2851] <= 3'b000;
      memory_array[2852] <= 3'b110;
      memory_array[2853] <= 3'b000;
      memory_array[2854] <= 3'b000;
      memory_array[2855] <= 3'b110;
      memory_array[2856] <= 3'b110;
      memory_array[2857] <= 3'b110;
      memory_array[2858] <= 3'b000;
      memory_array[2859] <= 3'b101;
      memory_array[2860] <= 3'b000;
      memory_array[2861] <= 3'b110;
      memory_array[2862] <= 3'b110;
      memory_array[2863] <= 3'b000;
      memory_array[2864] <= 3'b000;
      memory_array[2865] <= 3'b110;
      memory_array[2866] <= 3'b000;
      memory_array[2867] <= 3'b000;
      memory_array[2868] <= 3'b000;
      memory_array[2869] <= 3'b000;
      memory_array[2870] <= 3'b110;
      memory_array[2871] <= 3'b110;
      memory_array[2872] <= 3'b101;
      memory_array[2873] <= 3'b000;
      memory_array[2874] <= 3'b000;
      memory_array[2875] <= 3'b000;
      memory_array[2876] <= 3'b101;
      memory_array[2877] <= 3'b111;
      memory_array[2878] <= 3'b111;
      memory_array[2879] <= 3'b111;
      memory_array[2880] <= 3'b111;
      memory_array[2881] <= 3'b111;
      memory_array[2882] <= 3'b111;
      memory_array[2883] <= 3'b111;
      memory_array[2884] <= 3'b111;
      memory_array[2885] <= 3'b111;
      memory_array[2886] <= 3'b111;
      memory_array[2887] <= 3'b101;
      memory_array[2888] <= 3'b000;
      memory_array[2889] <= 3'b000;
      memory_array[2890] <= 3'b000;
      memory_array[2891] <= 3'b101;
      memory_array[2892] <= 3'b000;
      memory_array[2893] <= 3'b000;
      memory_array[2894] <= 3'b000;
      memory_array[2895] <= 3'b101;
      memory_array[2896] <= 3'b101;
      memory_array[2897] <= 3'b101;
      memory_array[2898] <= 3'b000;
      memory_array[2899] <= 3'b000;
      memory_array[2900] <= 3'b101;
      memory_array[2901] <= 3'b101;
      memory_array[2902] <= 3'b101;
      memory_array[2903] <= 3'b000;
      memory_array[2904] <= 3'b000;
      memory_array[2905] <= 3'b101;
      memory_array[2906] <= 3'b101;
      memory_array[2907] <= 3'b101;
      memory_array[2908] <= 3'b000;
      memory_array[2909] <= 3'b000;
      memory_array[2910] <= 3'b000;
      memory_array[2911] <= 3'b000;
      memory_array[2912] <= 3'b111;
      memory_array[2913] <= 3'b111;
      memory_array[2914] <= 3'b111;
      memory_array[2915] <= 3'b111;
      memory_array[2916] <= 3'b111;
      memory_array[2917] <= 3'b111;
      memory_array[2918] <= 3'b111;
      memory_array[2919] <= 3'b111;
      memory_array[2920] <= 3'b111;
      memory_array[2921] <= 3'b111;
      memory_array[2922] <= 3'b111;
      memory_array[2923] <= 3'b101;
      memory_array[2924] <= 3'b000;
      memory_array[2925] <= 3'b000;
      memory_array[2926] <= 3'b000;
      memory_array[2927] <= 3'b000;
      memory_array[2928] <= 3'b000;
      memory_array[2929] <= 3'b000;
      memory_array[2930] <= 3'b110;
      memory_array[2931] <= 3'b110;
      memory_array[2932] <= 3'b101;
      memory_array[2933] <= 3'b000;
      memory_array[2934] <= 3'b000;
      memory_array[2935] <= 3'b110;
      memory_array[2936] <= 3'b110;
      memory_array[2937] <= 3'b110;
      memory_array[2938] <= 3'b000;
      memory_array[2939] <= 3'b000;
      memory_array[2940] <= 3'b101;
      memory_array[2941] <= 3'b000;
      memory_array[2942] <= 3'b110;
      memory_array[2943] <= 3'b000;
      memory_array[2944] <= 3'b000;
      memory_array[2945] <= 3'b110;
      memory_array[2946] <= 3'b110;
      memory_array[2947] <= 3'b110;
      memory_array[2948] <= 3'b000;
      memory_array[2949] <= 3'b000;
      memory_array[2950] <= 3'b101;
      memory_array[2951] <= 3'b101;
      memory_array[2952] <= 3'b000;
      memory_array[2953] <= 3'b101;
      memory_array[2954] <= 3'b000;
      memory_array[2955] <= 3'b110;
      memory_array[2956] <= 3'b110;
      memory_array[2957] <= 3'b110;
      memory_array[2958] <= 3'b000;
      memory_array[2959] <= 3'b101;
      memory_array[2960] <= 3'b000;
      memory_array[2961] <= 3'b000;
      memory_array[2962] <= 3'b101;
      memory_array[2963] <= 3'b000;
      memory_array[2964] <= 3'b000;
      memory_array[2965] <= 3'b110;
      memory_array[2966] <= 3'b110;
      memory_array[2967] <= 3'b110;
      memory_array[2968] <= 3'b000;
      memory_array[2969] <= 3'b000;
      memory_array[2970] <= 3'b110;
      memory_array[2971] <= 3'b000;
      memory_array[2972] <= 3'b101;
      memory_array[2973] <= 3'b000;
      memory_array[2974] <= 3'b000;
      memory_array[2975] <= 3'b000;
      memory_array[2976] <= 3'b000;
      memory_array[2977] <= 3'b000;
      memory_array[2978] <= 3'b000;
      memory_array[2979] <= 3'b000;
      memory_array[2980] <= 3'b110;
      memory_array[2981] <= 3'b110;
      memory_array[2982] <= 3'b000;
      memory_array[2983] <= 3'b101;
      memory_array[2984] <= 3'b000;
      memory_array[2985] <= 3'b101;
      memory_array[2986] <= 3'b101;
      memory_array[2987] <= 3'b111;
      memory_array[2988] <= 3'b101;
      memory_array[2989] <= 3'b000;
      memory_array[2990] <= 3'b000;
      memory_array[2991] <= 3'b101;
      memory_array[2992] <= 3'b101;
      memory_array[2993] <= 3'b101;
      memory_array[2994] <= 3'b000;
      memory_array[2995] <= 3'b101;
      memory_array[2996] <= 3'b101;
      memory_array[2997] <= 3'b110;
      memory_array[2998] <= 3'b101;
      memory_array[2999] <= 3'b101;
      memory_array[3000] <= 3'b101;
      memory_array[3001] <= 3'b101;
      memory_array[3002] <= 3'b101;
      memory_array[3003] <= 3'b111;
      memory_array[3004] <= 3'b111;
      memory_array[3005] <= 3'b101;
      memory_array[3006] <= 3'b101;
      memory_array[3007] <= 3'b101;
      memory_array[3008] <= 3'b101;
      memory_array[3009] <= 3'b000;
      memory_array[3010] <= 3'b000;
      memory_array[3011] <= 3'b000;
      memory_array[3012] <= 3'b101;
      memory_array[3013] <= 3'b000;
      memory_array[3014] <= 3'b000;
      memory_array[3015] <= 3'b101;
      memory_array[3016] <= 3'b000;
      memory_array[3017] <= 3'b000;
      memory_array[3018] <= 3'b110;
      memory_array[3019] <= 3'b110;
      memory_array[3020] <= 3'b000;
      memory_array[3021] <= 3'b000;
      memory_array[3022] <= 3'b000;
      memory_array[3023] <= 3'b000;
      memory_array[3024] <= 3'b110;
      memory_array[3025] <= 3'b000;
      memory_array[3026] <= 3'b101;
      memory_array[3027] <= 3'b000;
      memory_array[3028] <= 3'b000;
      memory_array[3029] <= 3'b110;
      memory_array[3030] <= 3'b000;
      memory_array[3031] <= 3'b000;
      memory_array[3032] <= 3'b000;
      memory_array[3033] <= 3'b110;
      memory_array[3034] <= 3'b110;
      memory_array[3035] <= 3'b000;
      memory_array[3036] <= 3'b000;
      memory_array[3037] <= 3'b000;
      memory_array[3038] <= 3'b110;
      memory_array[3039] <= 3'b000;
      memory_array[3040] <= 3'b000;
      memory_array[3041] <= 3'b000;
      memory_array[3042] <= 3'b000;
      memory_array[3043] <= 3'b110;
      memory_array[3044] <= 3'b110;
      memory_array[3045] <= 3'b000;
      memory_array[3046] <= 3'b101;
      memory_array[3047] <= 3'b101;
      memory_array[3048] <= 3'b000;
      memory_array[3049] <= 3'b000;
      memory_array[3050] <= 3'b101;
      memory_array[3051] <= 3'b000;
      memory_array[3052] <= 3'b000;
      memory_array[3053] <= 3'b000;
      memory_array[3054] <= 3'b110;
      memory_array[3055] <= 3'b000;
      memory_array[3056] <= 3'b000;
      memory_array[3057] <= 3'b111;
      memory_array[3058] <= 3'b101;
      memory_array[3059] <= 3'b101;
      memory_array[3060] <= 3'b000;
      memory_array[3061] <= 3'b101;
      memory_array[3062] <= 3'b000;
      memory_array[3063] <= 3'b110;
      memory_array[3064] <= 3'b110;
      memory_array[3065] <= 3'b000;
      memory_array[3066] <= 3'b000;
      memory_array[3067] <= 3'b000;
      memory_array[3068] <= 3'b101;
      memory_array[3069] <= 3'b101;
      memory_array[3070] <= 3'b000;
      memory_array[3071] <= 3'b000;
      memory_array[3072] <= 3'b000;
      memory_array[3073] <= 3'b101;
      memory_array[3074] <= 3'b111;
      memory_array[3075] <= 3'b111;
      memory_array[3076] <= 3'b111;
      memory_array[3077] <= 3'b111;
      memory_array[3078] <= 3'b111;
      memory_array[3079] <= 3'b111;
      memory_array[3080] <= 3'b111;
      memory_array[3081] <= 3'b111;
      memory_array[3082] <= 3'b111;
      memory_array[3083] <= 3'b111;
      memory_array[3084] <= 3'b101;
      memory_array[3085] <= 3'b000;
      memory_array[3086] <= 3'b000;
      memory_array[3087] <= 3'b000;
      memory_array[3088] <= 3'b101;
      memory_array[3089] <= 3'b101;
      memory_array[3090] <= 3'b000;
      memory_array[3091] <= 3'b000;
      memory_array[3092] <= 3'b000;
      memory_array[3093] <= 3'b101;
      memory_array[3094] <= 3'b101;
      memory_array[3095] <= 3'b000;
      memory_array[3096] <= 3'b000;
      memory_array[3097] <= 3'b000;
      memory_array[3098] <= 3'b101;
      memory_array[3099] <= 3'b000;
      memory_array[3100] <= 3'b000;
      memory_array[3101] <= 3'b000;
      memory_array[3102] <= 3'b000;
      memory_array[3103] <= 3'b000;
      memory_array[3104] <= 3'b000;
      memory_array[3105] <= 3'b000;
      memory_array[3106] <= 3'b000;
      memory_array[3107] <= 3'b000;
      memory_array[3108] <= 3'b000;
      memory_array[3109] <= 3'b000;
      memory_array[3110] <= 3'b000;
      memory_array[3111] <= 3'b000;
      memory_array[3112] <= 3'b000;
      memory_array[3113] <= 3'b000;
      memory_array[3114] <= 3'b000;
      memory_array[3115] <= 3'b101;
      memory_array[3116] <= 3'b111;
      memory_array[3117] <= 3'b111;
      memory_array[3118] <= 3'b111;
      memory_array[3119] <= 3'b111;
      memory_array[3120] <= 3'b111;
      memory_array[3121] <= 3'b111;
      memory_array[3122] <= 3'b111;
      memory_array[3123] <= 3'b111;
      memory_array[3124] <= 3'b111;
      memory_array[3125] <= 3'b111;
      memory_array[3126] <= 3'b101;
      memory_array[3127] <= 3'b000;
      memory_array[3128] <= 3'b000;
      memory_array[3129] <= 3'b000;
      memory_array[3130] <= 3'b101;
      memory_array[3131] <= 3'b101;
      memory_array[3132] <= 3'b000;
      memory_array[3133] <= 3'b000;
      memory_array[3134] <= 3'b110;
      memory_array[3135] <= 3'b000;
      memory_array[3136] <= 3'b000;
      memory_array[3137] <= 3'b000;
      memory_array[3138] <= 3'b101;
      memory_array[3139] <= 3'b000;
      memory_array[3140] <= 3'b101;
      memory_array[3141] <= 3'b000;
      memory_array[3142] <= 3'b000;
      memory_array[3143] <= 3'b110;
      memory_array[3144] <= 3'b110;
      memory_array[3145] <= 3'b000;
      memory_array[3146] <= 3'b000;
      memory_array[3147] <= 3'b000;
      memory_array[3148] <= 3'b110;
      memory_array[3149] <= 3'b101;
      memory_array[3150] <= 3'b000;
      memory_array[3151] <= 3'b000;
      memory_array[3152] <= 3'b000;
      memory_array[3153] <= 3'b101;
      memory_array[3154] <= 3'b110;
      memory_array[3155] <= 3'b000;
      memory_array[3156] <= 3'b000;
      memory_array[3157] <= 3'b000;
      memory_array[3158] <= 3'b110;
      memory_array[3159] <= 3'b000;
      memory_array[3160] <= 3'b000;
      memory_array[3161] <= 3'b000;
      memory_array[3162] <= 3'b000;
      memory_array[3163] <= 3'b000;
      memory_array[3164] <= 3'b110;
      memory_array[3165] <= 3'b000;
      memory_array[3166] <= 3'b000;
      memory_array[3167] <= 3'b000;
      memory_array[3168] <= 3'b110;
      memory_array[3169] <= 3'b110;
      memory_array[3170] <= 3'b000;
      memory_array[3171] <= 3'b000;
      memory_array[3172] <= 3'b101;
      memory_array[3173] <= 3'b101;
      memory_array[3174] <= 3'b110;
      memory_array[3175] <= 3'b000;
      memory_array[3176] <= 3'b000;
      memory_array[3177] <= 3'b000;
      memory_array[3178] <= 3'b110;
      memory_array[3179] <= 3'b110;
      memory_array[3180] <= 3'b000;
      memory_array[3181] <= 3'b000;
      memory_array[3182] <= 3'b000;
      memory_array[3183] <= 3'b110;
      memory_array[3184] <= 3'b101;
      memory_array[3185] <= 3'b000;
      memory_array[3186] <= 3'b000;
      memory_array[3187] <= 3'b000;
      memory_array[3188] <= 3'b000;
      memory_array[3189] <= 3'b000;
      memory_array[3190] <= 3'b000;
      memory_array[3191] <= 3'b101;
      memory_array[3192] <= 3'b101;
      memory_array[3193] <= 3'b101;
      memory_array[3194] <= 3'b101;
      memory_array[3195] <= 3'b111;
      memory_array[3196] <= 3'b111;
      memory_array[3197] <= 3'b101;
      memory_array[3198] <= 3'b101;
      memory_array[3199] <= 3'b101;
      memory_array[3200] <= 3'b101;
      memory_array[3201] <= 3'b101;
      memory_array[3202] <= 3'b101;
      memory_array[3203] <= 3'b101;
      memory_array[3204] <= 3'b101;
      memory_array[3205] <= 3'b101;
      memory_array[3206] <= 3'b101;
      memory_array[3207] <= 3'b101;
      memory_array[3208] <= 3'b101;
      memory_array[3209] <= 3'b000;
      memory_array[3210] <= 3'b000;
      memory_array[3211] <= 3'b110;
      memory_array[3212] <= 3'b101;
      memory_array[3213] <= 3'b000;
      memory_array[3214] <= 3'b000;
      memory_array[3215] <= 3'b101;
      memory_array[3216] <= 3'b110;
      memory_array[3217] <= 3'b110;
      memory_array[3218] <= 3'b000;
      memory_array[3219] <= 3'b000;
      memory_array[3220] <= 3'b110;
      memory_array[3221] <= 3'b110;
      memory_array[3222] <= 3'b000;
      memory_array[3223] <= 3'b000;
      memory_array[3224] <= 3'b000;
      memory_array[3225] <= 3'b000;
      memory_array[3226] <= 3'b101;
      memory_array[3227] <= 3'b000;
      memory_array[3228] <= 3'b000;
      memory_array[3229] <= 3'b000;
      memory_array[3230] <= 3'b110;
      memory_array[3231] <= 3'b110;
      memory_array[3232] <= 3'b110;
      memory_array[3233] <= 3'b000;
      memory_array[3234] <= 3'b000;
      memory_array[3235] <= 3'b110;
      memory_array[3236] <= 3'b110;
      memory_array[3237] <= 3'b110;
      memory_array[3238] <= 3'b000;
      memory_array[3239] <= 3'b000;
      memory_array[3240] <= 3'b110;
      memory_array[3241] <= 3'b110;
      memory_array[3242] <= 3'b110;
      memory_array[3243] <= 3'b000;
      memory_array[3244] <= 3'b101;
      memory_array[3245] <= 3'b101;
      memory_array[3246] <= 3'b000;
      memory_array[3247] <= 3'b000;
      memory_array[3248] <= 3'b000;
      memory_array[3249] <= 3'b000;
      memory_array[3250] <= 3'b000;
      memory_array[3251] <= 3'b000;
      memory_array[3252] <= 3'b000;
      memory_array[3253] <= 3'b000;
      memory_array[3254] <= 3'b000;
      memory_array[3255] <= 3'b110;
      memory_array[3256] <= 3'b110;
      memory_array[3257] <= 3'b111;
      memory_array[3258] <= 3'b000;
      memory_array[3259] <= 3'b000;
      memory_array[3260] <= 3'b101;
      memory_array[3261] <= 3'b101;
      memory_array[3262] <= 3'b110;
      memory_array[3263] <= 3'b000;
      memory_array[3264] <= 3'b000;
      memory_array[3265] <= 3'b110;
      memory_array[3266] <= 3'b110;
      memory_array[3267] <= 3'b000;
      memory_array[3268] <= 3'b000;
      memory_array[3269] <= 3'b000;
      memory_array[3270] <= 3'b000;
      memory_array[3271] <= 3'b101;
      memory_array[3272] <= 3'b111;
      memory_array[3273] <= 3'b111;
      memory_array[3274] <= 3'b111;
      memory_array[3275] <= 3'b111;
      memory_array[3276] <= 3'b111;
      memory_array[3277] <= 3'b111;
      memory_array[3278] <= 3'b111;
      memory_array[3279] <= 3'b111;
      memory_array[3280] <= 3'b111;
      memory_array[3281] <= 3'b111;
      memory_array[3282] <= 3'b000;
      memory_array[3283] <= 3'b000;
      memory_array[3284] <= 3'b000;
      memory_array[3285] <= 3'b101;
      memory_array[3286] <= 3'b101;
      memory_array[3287] <= 3'b101;
      memory_array[3288] <= 3'b000;
      memory_array[3289] <= 3'b000;
      memory_array[3290] <= 3'b101;
      memory_array[3291] <= 3'b000;
      memory_array[3292] <= 3'b101;
      memory_array[3293] <= 3'b101;
      memory_array[3294] <= 3'b000;
      memory_array[3295] <= 3'b000;
      memory_array[3296] <= 3'b101;
      memory_array[3297] <= 3'b000;
      memory_array[3298] <= 3'b000;
      memory_array[3299] <= 3'b000;
      memory_array[3300] <= 3'b101;
      memory_array[3301] <= 3'b101;
      memory_array[3302] <= 3'b101;
      memory_array[3303] <= 3'b000;
      memory_array[3304] <= 3'b000;
      memory_array[3305] <= 3'b000;
      memory_array[3306] <= 3'b101;
      memory_array[3307] <= 3'b101;
      memory_array[3308] <= 3'b101;
      memory_array[3309] <= 3'b000;
      memory_array[3310] <= 3'b101;
      memory_array[3311] <= 3'b000;
      memory_array[3312] <= 3'b101;
      memory_array[3313] <= 3'b000;
      memory_array[3314] <= 3'b000;
      memory_array[3315] <= 3'b000;
      memory_array[3316] <= 3'b000;
      memory_array[3317] <= 3'b101;
      memory_array[3318] <= 3'b111;
      memory_array[3319] <= 3'b111;
      memory_array[3320] <= 3'b111;
      memory_array[3321] <= 3'b111;
      memory_array[3322] <= 3'b111;
      memory_array[3323] <= 3'b111;
      memory_array[3324] <= 3'b111;
      memory_array[3325] <= 3'b111;
      memory_array[3326] <= 3'b111;
      memory_array[3327] <= 3'b111;
      memory_array[3328] <= 3'b101;
      memory_array[3329] <= 3'b000;
      memory_array[3330] <= 3'b000;
      memory_array[3331] <= 3'b000;
      memory_array[3332] <= 3'b000;
      memory_array[3333] <= 3'b000;
      memory_array[3334] <= 3'b000;
      memory_array[3335] <= 3'b110;
      memory_array[3336] <= 3'b110;
      memory_array[3337] <= 3'b000;
      memory_array[3338] <= 3'b101;
      memory_array[3339] <= 3'b101;
      memory_array[3340] <= 3'b000;
      memory_array[3341] <= 3'b110;
      memory_array[3342] <= 3'b000;
      memory_array[3343] <= 3'b000;
      memory_array[3344] <= 3'b000;
      memory_array[3345] <= 3'b110;
      memory_array[3346] <= 3'b110;
      memory_array[3347] <= 3'b000;
      memory_array[3348] <= 3'b000;
      memory_array[3349] <= 3'b000;
      memory_array[3350] <= 3'b000;
      memory_array[3351] <= 3'b000;
      memory_array[3352] <= 3'b000;
      memory_array[3353] <= 3'b000;
      memory_array[3354] <= 3'b101;
      memory_array[3355] <= 3'b101;
      memory_array[3356] <= 3'b000;
      memory_array[3357] <= 3'b110;
      memory_array[3358] <= 3'b000;
      memory_array[3359] <= 3'b000;
      memory_array[3360] <= 3'b000;
      memory_array[3361] <= 3'b000;
      memory_array[3362] <= 3'b110;
      memory_array[3363] <= 3'b000;
      memory_array[3364] <= 3'b000;
      memory_array[3365] <= 3'b110;
      memory_array[3366] <= 3'b110;
      memory_array[3367] <= 3'b110;
      memory_array[3368] <= 3'b000;
      memory_array[3369] <= 3'b000;
      memory_array[3370] <= 3'b110;
      memory_array[3371] <= 3'b110;
      memory_array[3372] <= 3'b000;
      memory_array[3373] <= 3'b101;
      memory_array[3374] <= 3'b000;
      memory_array[3375] <= 3'b110;
      memory_array[3376] <= 3'b000;
      memory_array[3377] <= 3'b000;
      memory_array[3378] <= 3'b000;
      memory_array[3379] <= 3'b000;
      memory_array[3380] <= 3'b110;
      memory_array[3381] <= 3'b110;
      memory_array[3382] <= 3'b110;
      memory_array[3383] <= 3'b000;
      memory_array[3384] <= 3'b101;
      memory_array[3385] <= 3'b000;
      memory_array[3386] <= 3'b000;
      memory_array[3387] <= 3'b000;
      memory_array[3388] <= 3'b000;
      memory_array[3389] <= 3'b000;
      memory_array[3390] <= 3'b000;
      memory_array[3391] <= 3'b101;
      memory_array[3392] <= 3'b101;
      memory_array[3393] <= 3'b101;
      memory_array[3394] <= 3'b101;
      memory_array[3395] <= 3'b101;
      memory_array[3396] <= 3'b101;
      memory_array[3397] <= 3'b101;
      memory_array[3398] <= 3'b101;
      memory_array[3399] <= 3'b101;
      memory_array[3400] <= 3'b101;
      memory_array[3401] <= 3'b101;
      memory_array[3402] <= 3'b101;
      memory_array[3403] <= 3'b101;
      memory_array[3404] <= 3'b101;
      memory_array[3405] <= 3'b101;
      memory_array[3406] <= 3'b101;
      memory_array[3407] <= 3'b101;
      memory_array[3408] <= 3'b101;
      memory_array[3409] <= 3'b000;
      memory_array[3410] <= 3'b000;
      memory_array[3411] <= 3'b110;
      memory_array[3412] <= 3'b110;
      memory_array[3413] <= 3'b000;
      memory_array[3414] <= 3'b000;
      memory_array[3415] <= 3'b110;
      memory_array[3416] <= 3'b110;
      memory_array[3417] <= 3'b110;
      memory_array[3418] <= 3'b000;
      memory_array[3419] <= 3'b000;
      memory_array[3420] <= 3'b110;
      memory_array[3421] <= 3'b110;
      memory_array[3422] <= 3'b110;
      memory_array[3423] <= 3'b000;
      memory_array[3424] <= 3'b000;
      memory_array[3425] <= 3'b000;
      memory_array[3426] <= 3'b110;
      memory_array[3427] <= 3'b110;
      memory_array[3428] <= 3'b000;
      memory_array[3429] <= 3'b000;
      memory_array[3430] <= 3'b000;
      memory_array[3431] <= 3'b000;
      memory_array[3432] <= 3'b000;
      memory_array[3433] <= 3'b101;
      memory_array[3434] <= 3'b000;
      memory_array[3435] <= 3'b110;
      memory_array[3436] <= 3'b110;
      memory_array[3437] <= 3'b110;
      memory_array[3438] <= 3'b000;
      memory_array[3439] <= 3'b000;
      memory_array[3440] <= 3'b110;
      memory_array[3441] <= 3'b110;
      memory_array[3442] <= 3'b000;
      memory_array[3443] <= 3'b101;
      memory_array[3444] <= 3'b000;
      memory_array[3445] <= 3'b000;
      memory_array[3446] <= 3'b101;
      memory_array[3447] <= 3'b110;
      memory_array[3448] <= 3'b000;
      memory_array[3449] <= 3'b000;
      memory_array[3450] <= 3'b110;
      memory_array[3451] <= 3'b110;
      memory_array[3452] <= 3'b110;
      memory_array[3453] <= 3'b000;
      memory_array[3454] <= 3'b000;
      memory_array[3455] <= 3'b110;
      memory_array[3456] <= 3'b110;
      memory_array[3457] <= 3'b000;
      memory_array[3458] <= 3'b000;
      memory_array[3459] <= 3'b101;
      memory_array[3460] <= 3'b000;
      memory_array[3461] <= 3'b110;
      memory_array[3462] <= 3'b110;
      memory_array[3463] <= 3'b000;
      memory_array[3464] <= 3'b000;
      memory_array[3465] <= 3'b110;
      memory_array[3466] <= 3'b000;
      memory_array[3467] <= 3'b111;
      memory_array[3468] <= 3'b111;
      memory_array[3469] <= 3'b111;
      memory_array[3470] <= 3'b111;
      memory_array[3471] <= 3'b111;
      memory_array[3472] <= 3'b111;
      memory_array[3473] <= 3'b111;
      memory_array[3474] <= 3'b111;
      memory_array[3475] <= 3'b111;
      memory_array[3476] <= 3'b111;
      memory_array[3477] <= 3'b101;
      memory_array[3478] <= 3'b000;
      memory_array[3479] <= 3'b000;
      memory_array[3480] <= 3'b000;
      memory_array[3481] <= 3'b000;
      memory_array[3482] <= 3'b000;
      memory_array[3483] <= 3'b000;
      memory_array[3484] <= 3'b000;
      memory_array[3485] <= 3'b000;
      memory_array[3486] <= 3'b000;
      memory_array[3487] <= 3'b000;
      memory_array[3488] <= 3'b000;
      memory_array[3489] <= 3'b000;
      memory_array[3490] <= 3'b000;
      memory_array[3491] <= 3'b000;
      memory_array[3492] <= 3'b000;
      memory_array[3493] <= 3'b000;
      memory_array[3494] <= 3'b000;
      memory_array[3495] <= 3'b000;
      memory_array[3496] <= 3'b000;
      memory_array[3497] <= 3'b000;
      memory_array[3498] <= 3'b101;
      memory_array[3499] <= 3'b000;
      memory_array[3500] <= 3'b101;
      memory_array[3501] <= 3'b000;
      memory_array[3502] <= 3'b101;
      memory_array[3503] <= 3'b000;
      memory_array[3504] <= 3'b000;
      memory_array[3505] <= 3'b000;
      memory_array[3506] <= 3'b000;
      memory_array[3507] <= 3'b000;
      memory_array[3508] <= 3'b000;
      memory_array[3509] <= 3'b000;
      memory_array[3510] <= 3'b101;
      memory_array[3511] <= 3'b101;
      memory_array[3512] <= 3'b101;
      memory_array[3513] <= 3'b000;
      memory_array[3514] <= 3'b000;
      memory_array[3515] <= 3'b000;
      memory_array[3516] <= 3'b000;
      memory_array[3517] <= 3'b101;
      memory_array[3518] <= 3'b000;
      memory_array[3519] <= 3'b000;
      memory_array[3520] <= 3'b000;
      memory_array[3521] <= 3'b000;
      memory_array[3522] <= 3'b111;
      memory_array[3523] <= 3'b111;
      memory_array[3524] <= 3'b111;
      memory_array[3525] <= 3'b111;
      memory_array[3526] <= 3'b111;
      memory_array[3527] <= 3'b111;
      memory_array[3528] <= 3'b111;
      memory_array[3529] <= 3'b111;
      memory_array[3530] <= 3'b111;
      memory_array[3531] <= 3'b111;
      memory_array[3532] <= 3'b101;
      memory_array[3533] <= 3'b000;
      memory_array[3534] <= 3'b000;
      memory_array[3535] <= 3'b110;
      memory_array[3536] <= 3'b110;
      memory_array[3537] <= 3'b110;
      memory_array[3538] <= 3'b000;
      memory_array[3539] <= 3'b000;
      memory_array[3540] <= 3'b101;
      memory_array[3541] <= 3'b110;
      memory_array[3542] <= 3'b000;
      memory_array[3543] <= 3'b000;
      memory_array[3544] <= 3'b000;
      memory_array[3545] <= 3'b110;
      memory_array[3546] <= 3'b110;
      memory_array[3547] <= 3'b110;
      memory_array[3548] <= 3'b000;
      memory_array[3549] <= 3'b000;
      memory_array[3550] <= 3'b110;
      memory_array[3551] <= 3'b110;
      memory_array[3552] <= 3'b000;
      memory_array[3553] <= 3'b101;
      memory_array[3554] <= 3'b000;
      memory_array[3555] <= 3'b110;
      memory_array[3556] <= 3'b101;
      memory_array[3557] <= 3'b110;
      memory_array[3558] <= 3'b000;
      memory_array[3559] <= 3'b000;
      memory_array[3560] <= 3'b110;
      memory_array[3561] <= 3'b000;
      memory_array[3562] <= 3'b110;
      memory_array[3563] <= 3'b000;
      memory_array[3564] <= 3'b000;
      memory_array[3565] <= 3'b000;
      memory_array[3566] <= 3'b101;
      memory_array[3567] <= 3'b110;
      memory_array[3568] <= 3'b000;
      memory_array[3569] <= 3'b000;
      memory_array[3570] <= 3'b110;
      memory_array[3571] <= 3'b110;
      memory_array[3572] <= 3'b110;
      memory_array[3573] <= 3'b000;
      memory_array[3574] <= 3'b000;
      memory_array[3575] <= 3'b000;
      memory_array[3576] <= 3'b000;
      memory_array[3577] <= 3'b110;
      memory_array[3578] <= 3'b000;
      memory_array[3579] <= 3'b000;
      memory_array[3580] <= 3'b110;
      memory_array[3581] <= 3'b110;
      memory_array[3582] <= 3'b110;
      memory_array[3583] <= 3'b000;
      memory_array[3584] <= 3'b000;
      memory_array[3585] <= 3'b110;
      memory_array[3586] <= 3'b110;
      memory_array[3587] <= 3'b110;
      memory_array[3588] <= 3'b000;
      memory_array[3589] <= 3'b000;
      memory_array[3590] <= 3'b000;
      memory_array[3591] <= 3'b101;
      memory_array[3592] <= 3'b101;
      memory_array[3593] <= 3'b101;
      memory_array[3594] <= 3'b101;
      memory_array[3595] <= 3'b101;
      memory_array[3596] <= 3'b101;
      memory_array[3597] <= 3'b101;
      memory_array[3598] <= 3'b101;
      memory_array[3599] <= 3'b101;
      memory_array[3600] <= 3'b101;
      memory_array[3601] <= 3'b101;
      memory_array[3602] <= 3'b101;
      memory_array[3603] <= 3'b111;
      memory_array[3604] <= 3'b111;
      memory_array[3605] <= 3'b101;
      memory_array[3606] <= 3'b101;
      memory_array[3607] <= 3'b101;
      memory_array[3608] <= 3'b101;
      memory_array[3609] <= 3'b000;
      memory_array[3610] <= 3'b000;
      memory_array[3611] <= 3'b000;
      memory_array[3612] <= 3'b000;
      memory_array[3613] <= 3'b110;
      memory_array[3614] <= 3'b110;
      memory_array[3615] <= 3'b000;
      memory_array[3616] <= 3'b000;
      memory_array[3617] <= 3'b000;
      memory_array[3618] <= 3'b110;
      memory_array[3619] <= 3'b110;
      memory_array[3620] <= 3'b000;
      memory_array[3621] <= 3'b101;
      memory_array[3622] <= 3'b000;
      memory_array[3623] <= 3'b110;
      memory_array[3624] <= 3'b110;
      memory_array[3625] <= 3'b000;
      memory_array[3626] <= 3'b000;
      memory_array[3627] <= 3'b000;
      memory_array[3628] <= 3'b110;
      memory_array[3629] <= 3'b110;
      memory_array[3630] <= 3'b000;
      memory_array[3631] <= 3'b101;
      memory_array[3632] <= 3'b101;
      memory_array[3633] <= 3'b000;
      memory_array[3634] <= 3'b110;
      memory_array[3635] <= 3'b000;
      memory_array[3636] <= 3'b000;
      memory_array[3637] <= 3'b000;
      memory_array[3638] <= 3'b110;
      memory_array[3639] <= 3'b110;
      memory_array[3640] <= 3'b000;
      memory_array[3641] <= 3'b000;
      memory_array[3642] <= 3'b000;
      memory_array[3643] <= 3'b110;
      memory_array[3644] <= 3'b110;
      memory_array[3645] <= 3'b000;
      memory_array[3646] <= 3'b101;
      memory_array[3647] <= 3'b000;
      memory_array[3648] <= 3'b110;
      memory_array[3649] <= 3'b110;
      memory_array[3650] <= 3'b000;
      memory_array[3651] <= 3'b000;
      memory_array[3652] <= 3'b000;
      memory_array[3653] <= 3'b000;
      memory_array[3654] <= 3'b101;
      memory_array[3655] <= 3'b101;
      memory_array[3656] <= 3'b000;
      memory_array[3657] <= 3'b000;
      memory_array[3658] <= 3'b000;
      memory_array[3659] <= 3'b101;
      memory_array[3660] <= 3'b101;
      memory_array[3661] <= 3'b000;
      memory_array[3662] <= 3'b000;
      memory_array[3663] <= 3'b101;
      memory_array[3664] <= 3'b000;
      memory_array[3665] <= 3'b000;
      memory_array[3666] <= 3'b111;
      memory_array[3667] <= 3'b111;
      memory_array[3668] <= 3'b111;
      memory_array[3669] <= 3'b111;
      memory_array[3670] <= 3'b111;
      memory_array[3671] <= 3'b111;
      memory_array[3672] <= 3'b111;
      memory_array[3673] <= 3'b111;
      memory_array[3674] <= 3'b111;
      memory_array[3675] <= 3'b111;
      memory_array[3676] <= 3'b000;
      memory_array[3677] <= 3'b000;
      memory_array[3678] <= 3'b101;
      memory_array[3679] <= 3'b101;
      memory_array[3680] <= 3'b101;
      memory_array[3681] <= 3'b000;
      memory_array[3682] <= 3'b000;
      memory_array[3683] <= 3'b101;
      memory_array[3684] <= 3'b101;
      memory_array[3685] <= 3'b000;
      memory_array[3686] <= 3'b000;
      memory_array[3687] <= 3'b101;
      memory_array[3688] <= 3'b000;
      memory_array[3689] <= 3'b000;
      memory_array[3690] <= 3'b000;
      memory_array[3691] <= 3'b000;
      memory_array[3692] <= 3'b000;
      memory_array[3693] <= 3'b101;
      memory_array[3694] <= 3'b101;
      memory_array[3695] <= 3'b000;
      memory_array[3696] <= 3'b000;
      memory_array[3697] <= 3'b000;
      memory_array[3698] <= 3'b101;
      memory_array[3699] <= 3'b101;
      memory_array[3700] <= 3'b000;
      memory_array[3701] <= 3'b000;
      memory_array[3702] <= 3'b101;
      memory_array[3703] <= 3'b101;
      memory_array[3704] <= 3'b000;
      memory_array[3705] <= 3'b000;
      memory_array[3706] <= 3'b000;
      memory_array[3707] <= 3'b000;
      memory_array[3708] <= 3'b000;
      memory_array[3709] <= 3'b000;
      memory_array[3710] <= 3'b000;
      memory_array[3711] <= 3'b000;
      memory_array[3712] <= 3'b000;
      memory_array[3713] <= 3'b101;
      memory_array[3714] <= 3'b101;
      memory_array[3715] <= 3'b000;
      memory_array[3716] <= 3'b101;
      memory_array[3717] <= 3'b000;
      memory_array[3718] <= 3'b101;
      memory_array[3719] <= 3'b101;
      memory_array[3720] <= 3'b000;
      memory_array[3721] <= 3'b000;
      memory_array[3722] <= 3'b000;
      memory_array[3723] <= 3'b000;
      memory_array[3724] <= 3'b111;
      memory_array[3725] <= 3'b111;
      memory_array[3726] <= 3'b111;
      memory_array[3727] <= 3'b111;
      memory_array[3728] <= 3'b111;
      memory_array[3729] <= 3'b111;
      memory_array[3730] <= 3'b111;
      memory_array[3731] <= 3'b111;
      memory_array[3732] <= 3'b111;
      memory_array[3733] <= 3'b111;
      memory_array[3734] <= 3'b000;
      memory_array[3735] <= 3'b000;
      memory_array[3736] <= 3'b000;
      memory_array[3737] <= 3'b000;
      memory_array[3738] <= 3'b110;
      memory_array[3739] <= 3'b101;
      memory_array[3740] <= 3'b101;
      memory_array[3741] <= 3'b000;
      memory_array[3742] <= 3'b000;
      memory_array[3743] <= 3'b000;
      memory_array[3744] <= 3'b101;
      memory_array[3745] <= 3'b101;
      memory_array[3746] <= 3'b000;
      memory_array[3747] <= 3'b000;
      memory_array[3748] <= 3'b110;
      memory_array[3749] <= 3'b110;
      memory_array[3750] <= 3'b000;
      memory_array[3751] <= 3'b000;
      memory_array[3752] <= 3'b000;
      memory_array[3753] <= 3'b101;
      memory_array[3754] <= 3'b110;
      memory_array[3755] <= 3'b000;
      memory_array[3756] <= 3'b000;
      memory_array[3757] <= 3'b000;
      memory_array[3758] <= 3'b110;
      memory_array[3759] <= 3'b110;
      memory_array[3760] <= 3'b000;
      memory_array[3761] <= 3'b000;
      memory_array[3762] <= 3'b000;
      memory_array[3763] <= 3'b110;
      memory_array[3764] <= 3'b110;
      memory_array[3765] <= 3'b000;
      memory_array[3766] <= 3'b000;
      memory_array[3767] <= 3'b101;
      memory_array[3768] <= 3'b101;
      memory_array[3769] <= 3'b000;
      memory_array[3770] <= 3'b000;
      memory_array[3771] <= 3'b000;
      memory_array[3772] <= 3'b000;
      memory_array[3773] <= 3'b000;
      memory_array[3774] <= 3'b000;
      memory_array[3775] <= 3'b000;
      memory_array[3776] <= 3'b000;
      memory_array[3777] <= 3'b101;
      memory_array[3778] <= 3'b101;
      memory_array[3779] <= 3'b110;
      memory_array[3780] <= 3'b000;
      memory_array[3781] <= 3'b000;
      memory_array[3782] <= 3'b000;
      memory_array[3783] <= 3'b110;
      memory_array[3784] <= 3'b110;
      memory_array[3785] <= 3'b000;
      memory_array[3786] <= 3'b000;
      memory_array[3787] <= 3'b000;
      memory_array[3788] <= 3'b110;
      memory_array[3789] <= 3'b000;
      memory_array[3790] <= 3'b000;
      memory_array[3791] <= 3'b101;
      memory_array[3792] <= 3'b101;
      memory_array[3793] <= 3'b101;
      memory_array[3794] <= 3'b101;
      memory_array[3795] <= 3'b111;
      memory_array[3796] <= 3'b111;
      memory_array[3797] <= 3'b101;
      memory_array[3798] <= 3'b101;
      memory_array[3799] <= 3'b101;
      memory_array[3800] <= 3'b101;
      memory_array[3801] <= 3'b000;
      memory_array[3802] <= 3'b000;
      memory_array[3803] <= 3'b110;
      memory_array[3804] <= 3'b110;
      memory_array[3805] <= 3'b000;
      memory_array[3806] <= 3'b000;
      memory_array[3807] <= 3'b101;
      memory_array[3808] <= 3'b101;
      memory_array[3809] <= 3'b000;
      memory_array[3810] <= 3'b000;
      memory_array[3811] <= 3'b000;
      memory_array[3812] <= 3'b000;
      memory_array[3813] <= 3'b110;
      memory_array[3814] <= 3'b110;
      memory_array[3815] <= 3'b000;
      memory_array[3816] <= 3'b000;
      memory_array[3817] <= 3'b000;
      memory_array[3818] <= 3'b110;
      memory_array[3819] <= 3'b110;
      memory_array[3820] <= 3'b000;
      memory_array[3821] <= 3'b000;
      memory_array[3822] <= 3'b000;
      memory_array[3823] <= 3'b110;
      memory_array[3824] <= 3'b110;
      memory_array[3825] <= 3'b000;
      memory_array[3826] <= 3'b000;
      memory_array[3827] <= 3'b101;
      memory_array[3828] <= 3'b101;
      memory_array[3829] <= 3'b000;
      memory_array[3830] <= 3'b000;
      memory_array[3831] <= 3'b101;
      memory_array[3832] <= 3'b000;
      memory_array[3833] <= 3'b110;
      memory_array[3834] <= 3'b110;
      memory_array[3835] <= 3'b000;
      memory_array[3836] <= 3'b000;
      memory_array[3837] <= 3'b000;
      memory_array[3838] <= 3'b110;
      memory_array[3839] <= 3'b110;
      memory_array[3840] <= 3'b000;
      memory_array[3841] <= 3'b000;
      memory_array[3842] <= 3'b000;
      memory_array[3843] <= 3'b110;
      memory_array[3844] <= 3'b110;
      memory_array[3845] <= 3'b000;
      memory_array[3846] <= 3'b000;
      memory_array[3847] <= 3'b000;
      memory_array[3848] <= 3'b110;
      memory_array[3849] <= 3'b110;
      memory_array[3850] <= 3'b000;
      memory_array[3851] <= 3'b000;
      memory_array[3852] <= 3'b000;
      memory_array[3853] <= 3'b101;
      memory_array[3854] <= 3'b000;
      memory_array[3855] <= 3'b000;
      memory_array[3856] <= 3'b101;
      memory_array[3857] <= 3'b000;
      memory_array[3858] <= 3'b101;
      memory_array[3859] <= 3'b000;
      memory_array[3860] <= 3'b000;
      memory_array[3861] <= 3'b000;
      memory_array[3862] <= 3'b101;
      memory_array[3863] <= 3'b111;
      memory_array[3864] <= 3'b111;
      memory_array[3865] <= 3'b111;
      memory_array[3866] <= 3'b111;
      memory_array[3867] <= 3'b111;
      memory_array[3868] <= 3'b111;
      memory_array[3869] <= 3'b111;
      memory_array[3870] <= 3'b111;
      memory_array[3871] <= 3'b111;
      memory_array[3872] <= 3'b000;
      memory_array[3873] <= 3'b000;
      memory_array[3874] <= 3'b101;
      memory_array[3875] <= 3'b000;
      memory_array[3876] <= 3'b000;
      memory_array[3877] <= 3'b000;
      memory_array[3878] <= 3'b000;
      memory_array[3879] <= 3'b101;
      memory_array[3880] <= 3'b000;
      memory_array[3881] <= 3'b000;
      memory_array[3882] <= 3'b101;
      memory_array[3883] <= 3'b101;
      memory_array[3884] <= 3'b000;
      memory_array[3885] <= 3'b000;
      memory_array[3886] <= 3'b000;
      memory_array[3887] <= 3'b101;
      memory_array[3888] <= 3'b000;
      memory_array[3889] <= 3'b000;
      memory_array[3890] <= 3'b000;
      memory_array[3891] <= 3'b000;
      memory_array[3892] <= 3'b000;
      memory_array[3893] <= 3'b101;
      memory_array[3894] <= 3'b101;
      memory_array[3895] <= 3'b101;
      memory_array[3896] <= 3'b000;
      memory_array[3897] <= 3'b000;
      memory_array[3898] <= 3'b101;
      memory_array[3899] <= 3'b101;
      memory_array[3900] <= 3'b101;
      memory_array[3901] <= 3'b101;
      memory_array[3902] <= 3'b000;
      memory_array[3903] <= 3'b000;
      memory_array[3904] <= 3'b101;
      memory_array[3905] <= 3'b000;
      memory_array[3906] <= 3'b000;
      memory_array[3907] <= 3'b000;
      memory_array[3908] <= 3'b101;
      memory_array[3909] <= 3'b101;
      memory_array[3910] <= 3'b101;
      memory_array[3911] <= 3'b000;
      memory_array[3912] <= 3'b000;
      memory_array[3913] <= 3'b101;
      memory_array[3914] <= 3'b101;
      memory_array[3915] <= 3'b000;
      memory_array[3916] <= 3'b000;
      memory_array[3917] <= 3'b000;
      memory_array[3918] <= 3'b101;
      memory_array[3919] <= 3'b000;
      memory_array[3920] <= 3'b101;
      memory_array[3921] <= 3'b000;
      memory_array[3922] <= 3'b000;
      memory_array[3923] <= 3'b000;
      memory_array[3924] <= 3'b101;
      memory_array[3925] <= 3'b000;
      memory_array[3926] <= 3'b000;
      memory_array[3927] <= 3'b101;
      memory_array[3928] <= 3'b111;
      memory_array[3929] <= 3'b111;
      memory_array[3930] <= 3'b111;
      memory_array[3931] <= 3'b111;
      memory_array[3932] <= 3'b111;
      memory_array[3933] <= 3'b111;
      memory_array[3934] <= 3'b111;
      memory_array[3935] <= 3'b111;
      memory_array[3936] <= 3'b111;
      memory_array[3937] <= 3'b000;
      memory_array[3938] <= 3'b000;
      memory_array[3939] <= 3'b000;
      memory_array[3940] <= 3'b000;
      memory_array[3941] <= 3'b101;
      memory_array[3942] <= 3'b000;
      memory_array[3943] <= 3'b101;
      memory_array[3944] <= 3'b000;
      memory_array[3945] <= 3'b000;
      memory_array[3946] <= 3'b101;
      memory_array[3947] <= 3'b000;
      memory_array[3948] <= 3'b110;
      memory_array[3949] <= 3'b110;
      memory_array[3950] <= 3'b000;
      memory_array[3951] <= 3'b000;
      memory_array[3952] <= 3'b101;
      memory_array[3953] <= 3'b000;
      memory_array[3954] <= 3'b110;
      memory_array[3955] <= 3'b000;
      memory_array[3956] <= 3'b000;
      memory_array[3957] <= 3'b000;
      memory_array[3958] <= 3'b110;
      memory_array[3959] <= 3'b110;
      memory_array[3960] <= 3'b000;
      memory_array[3961] <= 3'b000;
      memory_array[3962] <= 3'b000;
      memory_array[3963] <= 3'b110;
      memory_array[3964] <= 3'b110;
      memory_array[3965] <= 3'b000;
      memory_array[3966] <= 3'b000;
      memory_array[3967] <= 3'b000;
      memory_array[3968] <= 3'b101;
      memory_array[3969] <= 3'b000;
      memory_array[3970] <= 3'b000;
      memory_array[3971] <= 3'b101;
      memory_array[3972] <= 3'b101;
      memory_array[3973] <= 3'b000;
      memory_array[3974] <= 3'b110;
      memory_array[3975] <= 3'b000;
      memory_array[3976] <= 3'b000;
      memory_array[3977] <= 3'b000;
      memory_array[3978] <= 3'b000;
      memory_array[3979] <= 3'b110;
      memory_array[3980] <= 3'b000;
      memory_array[3981] <= 3'b000;
      memory_array[3982] <= 3'b000;
      memory_array[3983] <= 3'b110;
      memory_array[3984] <= 3'b110;
      memory_array[3985] <= 3'b000;
      memory_array[3986] <= 3'b000;
      memory_array[3987] <= 3'b000;
      memory_array[3988] <= 3'b110;
      memory_array[3989] <= 3'b000;
      memory_array[3990] <= 3'b000;
      memory_array[3991] <= 3'b101;
      memory_array[3992] <= 3'b101;
      memory_array[3993] <= 3'b110;
      memory_array[3994] <= 3'b110;
      memory_array[3995] <= 3'b000;
      memory_array[3996] <= 3'b000;
      memory_array[3997] <= 3'b000;
      memory_array[3998] <= 3'b110;
      memory_array[3999] <= 3'b101;
      memory_array[4000] <= 3'b101;
      memory_array[4001] <= 3'b000;
      memory_array[4002] <= 3'b000;
      memory_array[4003] <= 3'b110;
      memory_array[4004] <= 3'b110;
      memory_array[4005] <= 3'b000;
      memory_array[4006] <= 3'b000;
      memory_array[4007] <= 3'b101;
      memory_array[4008] <= 3'b101;
      memory_array[4009] <= 3'b000;
      memory_array[4010] <= 3'b000;
      memory_array[4011] <= 3'b000;
      memory_array[4012] <= 3'b000;
      memory_array[4013] <= 3'b110;
      memory_array[4014] <= 3'b110;
      memory_array[4015] <= 3'b000;
      memory_array[4016] <= 3'b000;
      memory_array[4017] <= 3'b000;
      memory_array[4018] <= 3'b110;
      memory_array[4019] <= 3'b110;
      memory_array[4020] <= 3'b000;
      memory_array[4021] <= 3'b000;
      memory_array[4022] <= 3'b000;
      memory_array[4023] <= 3'b110;
      memory_array[4024] <= 3'b110;
      memory_array[4025] <= 3'b000;
      memory_array[4026] <= 3'b000;
      memory_array[4027] <= 3'b101;
      memory_array[4028] <= 3'b101;
      memory_array[4029] <= 3'b000;
      memory_array[4030] <= 3'b000;
      memory_array[4031] <= 3'b101;
      memory_array[4032] <= 3'b000;
      memory_array[4033] <= 3'b110;
      memory_array[4034] <= 3'b110;
      memory_array[4035] <= 3'b000;
      memory_array[4036] <= 3'b000;
      memory_array[4037] <= 3'b000;
      memory_array[4038] <= 3'b110;
      memory_array[4039] <= 3'b110;
      memory_array[4040] <= 3'b000;
      memory_array[4041] <= 3'b000;
      memory_array[4042] <= 3'b000;
      memory_array[4043] <= 3'b110;
      memory_array[4044] <= 3'b110;
      memory_array[4045] <= 3'b000;
      memory_array[4046] <= 3'b000;
      memory_array[4047] <= 3'b000;
      memory_array[4048] <= 3'b110;
      memory_array[4049] <= 3'b110;
      memory_array[4050] <= 3'b000;
      memory_array[4051] <= 3'b000;
      memory_array[4052] <= 3'b000;
      memory_array[4053] <= 3'b101;
      memory_array[4054] <= 3'b000;
      memory_array[4055] <= 3'b000;
      memory_array[4056] <= 3'b101;
      memory_array[4057] <= 3'b000;
      memory_array[4058] <= 3'b101;
      memory_array[4059] <= 3'b000;
      memory_array[4060] <= 3'b000;
      memory_array[4061] <= 3'b000;
      memory_array[4062] <= 3'b101;
      memory_array[4063] <= 3'b111;
      memory_array[4064] <= 3'b111;
      memory_array[4065] <= 3'b111;
      memory_array[4066] <= 3'b111;
      memory_array[4067] <= 3'b111;
      memory_array[4068] <= 3'b111;
      memory_array[4069] <= 3'b111;
      memory_array[4070] <= 3'b111;
      memory_array[4071] <= 3'b111;
      memory_array[4072] <= 3'b000;
      memory_array[4073] <= 3'b000;
      memory_array[4074] <= 3'b101;
      memory_array[4075] <= 3'b000;
      memory_array[4076] <= 3'b000;
      memory_array[4077] <= 3'b000;
      memory_array[4078] <= 3'b000;
      memory_array[4079] <= 3'b101;
      memory_array[4080] <= 3'b000;
      memory_array[4081] <= 3'b000;
      memory_array[4082] <= 3'b101;
      memory_array[4083] <= 3'b101;
      memory_array[4084] <= 3'b000;
      memory_array[4085] <= 3'b000;
      memory_array[4086] <= 3'b000;
      memory_array[4087] <= 3'b101;
      memory_array[4088] <= 3'b000;
      memory_array[4089] <= 3'b000;
      memory_array[4090] <= 3'b000;
      memory_array[4091] <= 3'b000;
      memory_array[4092] <= 3'b000;
      memory_array[4093] <= 3'b101;
      memory_array[4094] <= 3'b101;
      memory_array[4095] <= 3'b101;
      memory_array[4096] <= 3'b000;
      memory_array[4097] <= 3'b000;
      memory_array[4098] <= 3'b101;
      memory_array[4099] <= 3'b101;
      memory_array[4100] <= 3'b101;
      memory_array[4101] <= 3'b101;
      memory_array[4102] <= 3'b000;
      memory_array[4103] <= 3'b000;
      memory_array[4104] <= 3'b101;
      memory_array[4105] <= 3'b000;
      memory_array[4106] <= 3'b000;
      memory_array[4107] <= 3'b000;
      memory_array[4108] <= 3'b101;
      memory_array[4109] <= 3'b101;
      memory_array[4110] <= 3'b101;
      memory_array[4111] <= 3'b000;
      memory_array[4112] <= 3'b000;
      memory_array[4113] <= 3'b101;
      memory_array[4114] <= 3'b101;
      memory_array[4115] <= 3'b000;
      memory_array[4116] <= 3'b000;
      memory_array[4117] <= 3'b000;
      memory_array[4118] <= 3'b101;
      memory_array[4119] <= 3'b000;
      memory_array[4120] <= 3'b101;
      memory_array[4121] <= 3'b000;
      memory_array[4122] <= 3'b000;
      memory_array[4123] <= 3'b000;
      memory_array[4124] <= 3'b101;
      memory_array[4125] <= 3'b000;
      memory_array[4126] <= 3'b000;
      memory_array[4127] <= 3'b101;
      memory_array[4128] <= 3'b111;
      memory_array[4129] <= 3'b111;
      memory_array[4130] <= 3'b111;
      memory_array[4131] <= 3'b111;
      memory_array[4132] <= 3'b111;
      memory_array[4133] <= 3'b111;
      memory_array[4134] <= 3'b111;
      memory_array[4135] <= 3'b111;
      memory_array[4136] <= 3'b111;
      memory_array[4137] <= 3'b000;
      memory_array[4138] <= 3'b000;
      memory_array[4139] <= 3'b000;
      memory_array[4140] <= 3'b000;
      memory_array[4141] <= 3'b101;
      memory_array[4142] <= 3'b000;
      memory_array[4143] <= 3'b101;
      memory_array[4144] <= 3'b000;
      memory_array[4145] <= 3'b000;
      memory_array[4146] <= 3'b101;
      memory_array[4147] <= 3'b000;
      memory_array[4148] <= 3'b110;
      memory_array[4149] <= 3'b110;
      memory_array[4150] <= 3'b000;
      memory_array[4151] <= 3'b000;
      memory_array[4152] <= 3'b101;
      memory_array[4153] <= 3'b000;
      memory_array[4154] <= 3'b110;
      memory_array[4155] <= 3'b000;
      memory_array[4156] <= 3'b000;
      memory_array[4157] <= 3'b000;
      memory_array[4158] <= 3'b110;
      memory_array[4159] <= 3'b110;
      memory_array[4160] <= 3'b000;
      memory_array[4161] <= 3'b000;
      memory_array[4162] <= 3'b000;
      memory_array[4163] <= 3'b110;
      memory_array[4164] <= 3'b110;
      memory_array[4165] <= 3'b000;
      memory_array[4166] <= 3'b000;
      memory_array[4167] <= 3'b000;
      memory_array[4168] <= 3'b101;
      memory_array[4169] <= 3'b000;
      memory_array[4170] <= 3'b000;
      memory_array[4171] <= 3'b101;
      memory_array[4172] <= 3'b101;
      memory_array[4173] <= 3'b000;
      memory_array[4174] <= 3'b110;
      memory_array[4175] <= 3'b000;
      memory_array[4176] <= 3'b000;
      memory_array[4177] <= 3'b000;
      memory_array[4178] <= 3'b000;
      memory_array[4179] <= 3'b110;
      memory_array[4180] <= 3'b000;
      memory_array[4181] <= 3'b000;
      memory_array[4182] <= 3'b000;
      memory_array[4183] <= 3'b110;
      memory_array[4184] <= 3'b110;
      memory_array[4185] <= 3'b000;
      memory_array[4186] <= 3'b000;
      memory_array[4187] <= 3'b000;
      memory_array[4188] <= 3'b110;
      memory_array[4189] <= 3'b000;
      memory_array[4190] <= 3'b000;
      memory_array[4191] <= 3'b101;
      memory_array[4192] <= 3'b101;
      memory_array[4193] <= 3'b110;
      memory_array[4194] <= 3'b110;
      memory_array[4195] <= 3'b000;
      memory_array[4196] <= 3'b000;
      memory_array[4197] <= 3'b000;
      memory_array[4198] <= 3'b110;
      memory_array[4199] <= 3'b101;
      memory_array[4200] <= 3'b000;
      memory_array[4201] <= 3'b000;
      memory_array[4202] <= 3'b000;
      memory_array[4203] <= 3'b110;
      memory_array[4204] <= 3'b110;
      memory_array[4205] <= 3'b000;
      memory_array[4206] <= 3'b000;
      memory_array[4207] <= 3'b000;
      memory_array[4208] <= 3'b101;
      memory_array[4209] <= 3'b000;
      memory_array[4210] <= 3'b000;
      memory_array[4211] <= 3'b000;
      memory_array[4212] <= 3'b000;
      memory_array[4213] <= 3'b110;
      memory_array[4214] <= 3'b110;
      memory_array[4215] <= 3'b000;
      memory_array[4216] <= 3'b000;
      memory_array[4217] <= 3'b000;
      memory_array[4218] <= 3'b101;
      memory_array[4219] <= 3'b110;
      memory_array[4220] <= 3'b000;
      memory_array[4221] <= 3'b000;
      memory_array[4222] <= 3'b000;
      memory_array[4223] <= 3'b000;
      memory_array[4224] <= 3'b101;
      memory_array[4225] <= 3'b000;
      memory_array[4226] <= 3'b000;
      memory_array[4227] <= 3'b000;
      memory_array[4228] <= 3'b000;
      memory_array[4229] <= 3'b000;
      memory_array[4230] <= 3'b000;
      memory_array[4231] <= 3'b000;
      memory_array[4232] <= 3'b000;
      memory_array[4233] <= 3'b110;
      memory_array[4234] <= 3'b110;
      memory_array[4235] <= 3'b000;
      memory_array[4236] <= 3'b000;
      memory_array[4237] <= 3'b000;
      memory_array[4238] <= 3'b110;
      memory_array[4239] <= 3'b110;
      memory_array[4240] <= 3'b000;
      memory_array[4241] <= 3'b000;
      memory_array[4242] <= 3'b000;
      memory_array[4243] <= 3'b110;
      memory_array[4244] <= 3'b110;
      memory_array[4245] <= 3'b000;
      memory_array[4246] <= 3'b000;
      memory_array[4247] <= 3'b000;
      memory_array[4248] <= 3'b101;
      memory_array[4249] <= 3'b110;
      memory_array[4250] <= 3'b000;
      memory_array[4251] <= 3'b000;
      memory_array[4252] <= 3'b000;
      memory_array[4253] <= 3'b110;
      memory_array[4254] <= 3'b110;
      memory_array[4255] <= 3'b000;
      memory_array[4256] <= 3'b101;
      memory_array[4257] <= 3'b000;
      memory_array[4258] <= 3'b000;
      memory_array[4259] <= 3'b101;
      memory_array[4260] <= 3'b111;
      memory_array[4261] <= 3'b111;
      memory_array[4262] <= 3'b111;
      memory_array[4263] <= 3'b111;
      memory_array[4264] <= 3'b111;
      memory_array[4265] <= 3'b111;
      memory_array[4266] <= 3'b111;
      memory_array[4267] <= 3'b111;
      memory_array[4268] <= 3'b101;
      memory_array[4269] <= 3'b000;
      memory_array[4270] <= 3'b000;
      memory_array[4271] <= 3'b000;
      memory_array[4272] <= 3'b101;
      memory_array[4273] <= 3'b000;
      memory_array[4274] <= 3'b101;
      memory_array[4275] <= 3'b000;
      memory_array[4276] <= 3'b000;
      memory_array[4277] <= 3'b000;
      memory_array[4278] <= 3'b101;
      memory_array[4279] <= 3'b101;
      memory_array[4280] <= 3'b000;
      memory_array[4281] <= 3'b101;
      memory_array[4282] <= 3'b000;
      memory_array[4283] <= 3'b000;
      memory_array[4284] <= 3'b101;
      memory_array[4285] <= 3'b000;
      memory_array[4286] <= 3'b000;
      memory_array[4287] <= 3'b000;
      memory_array[4288] <= 3'b000;
      memory_array[4289] <= 3'b101;
      memory_array[4290] <= 3'b000;
      memory_array[4291] <= 3'b101;
      memory_array[4292] <= 3'b000;
      memory_array[4293] <= 3'b000;
      memory_array[4294] <= 3'b101;
      memory_array[4295] <= 3'b000;
      memory_array[4296] <= 3'b000;
      memory_array[4297] <= 3'b101;
      memory_array[4298] <= 3'b101;
      memory_array[4299] <= 3'b101;
      memory_array[4300] <= 3'b000;
      memory_array[4301] <= 3'b000;
      memory_array[4302] <= 3'b000;
      memory_array[4303] <= 3'b000;
      memory_array[4304] <= 3'b101;
      memory_array[4305] <= 3'b000;
      memory_array[4306] <= 3'b000;
      memory_array[4307] <= 3'b101;
      memory_array[4308] <= 3'b000;
      memory_array[4309] <= 3'b101;
      memory_array[4310] <= 3'b000;
      memory_array[4311] <= 3'b000;
      memory_array[4312] <= 3'b000;
      memory_array[4313] <= 3'b101;
      memory_array[4314] <= 3'b000;
      memory_array[4315] <= 3'b000;
      memory_array[4316] <= 3'b000;
      memory_array[4317] <= 3'b000;
      memory_array[4318] <= 3'b101;
      memory_array[4319] <= 3'b101;
      memory_array[4320] <= 3'b000;
      memory_array[4321] <= 3'b000;
      memory_array[4322] <= 3'b000;
      memory_array[4323] <= 3'b000;
      memory_array[4324] <= 3'b101;
      memory_array[4325] <= 3'b000;
      memory_array[4326] <= 3'b000;
      memory_array[4327] <= 3'b101;
      memory_array[4328] <= 3'b000;
      memory_array[4329] <= 3'b000;
      memory_array[4330] <= 3'b000;
      memory_array[4331] <= 3'b101;
      memory_array[4332] <= 3'b111;
      memory_array[4333] <= 3'b111;
      memory_array[4334] <= 3'b111;
      memory_array[4335] <= 3'b111;
      memory_array[4336] <= 3'b111;
      memory_array[4337] <= 3'b111;
      memory_array[4338] <= 3'b111;
      memory_array[4339] <= 3'b111;
      memory_array[4340] <= 3'b101;
      memory_array[4341] <= 3'b000;
      memory_array[4342] <= 3'b000;
      memory_array[4343] <= 3'b101;
      memory_array[4344] <= 3'b110;
      memory_array[4345] <= 3'b000;
      memory_array[4346] <= 3'b000;
      memory_array[4347] <= 3'b000;
      memory_array[4348] <= 3'b110;
      memory_array[4349] <= 3'b110;
      memory_array[4350] <= 3'b000;
      memory_array[4351] <= 3'b101;
      memory_array[4352] <= 3'b000;
      memory_array[4353] <= 3'b000;
      memory_array[4354] <= 3'b000;
      memory_array[4355] <= 3'b000;
      memory_array[4356] <= 3'b000;
      memory_array[4357] <= 3'b000;
      memory_array[4358] <= 3'b110;
      memory_array[4359] <= 3'b110;
      memory_array[4360] <= 3'b000;
      memory_array[4361] <= 3'b000;
      memory_array[4362] <= 3'b000;
      memory_array[4363] <= 3'b110;
      memory_array[4364] <= 3'b110;
      memory_array[4365] <= 3'b000;
      memory_array[4366] <= 3'b000;
      memory_array[4367] <= 3'b000;
      memory_array[4368] <= 3'b110;
      memory_array[4369] <= 3'b000;
      memory_array[4370] <= 3'b000;
      memory_array[4371] <= 3'b000;
      memory_array[4372] <= 3'b000;
      memory_array[4373] <= 3'b000;
      memory_array[4374] <= 3'b000;
      memory_array[4375] <= 3'b101;
      memory_array[4376] <= 3'b000;
      memory_array[4377] <= 3'b000;
      memory_array[4378] <= 3'b110;
      memory_array[4379] <= 3'b110;
      memory_array[4380] <= 3'b000;
      memory_array[4381] <= 3'b101;
      memory_array[4382] <= 3'b000;
      memory_array[4383] <= 3'b110;
      memory_array[4384] <= 3'b110;
      memory_array[4385] <= 3'b000;
      memory_array[4386] <= 3'b000;
      memory_array[4387] <= 3'b000;
      memory_array[4388] <= 3'b110;
      memory_array[4389] <= 3'b000;
      memory_array[4390] <= 3'b000;
      memory_array[4391] <= 3'b101;
      memory_array[4392] <= 3'b000;
      memory_array[4393] <= 3'b110;
      memory_array[4394] <= 3'b110;
      memory_array[4395] <= 3'b000;
      memory_array[4396] <= 3'b000;
      memory_array[4397] <= 3'b000;
      memory_array[4398] <= 3'b110;
      memory_array[4399] <= 3'b110;
      memory_array[4400] <= 3'b101;
      memory_array[4401] <= 3'b101;
      memory_array[4402] <= 3'b101;
      memory_array[4403] <= 3'b101;
      memory_array[4404] <= 3'b101;
      memory_array[4405] <= 3'b101;
      memory_array[4406] <= 3'b101;
      memory_array[4407] <= 3'b101;
      memory_array[4408] <= 3'b101;
      memory_array[4409] <= 3'b000;
      memory_array[4410] <= 3'b000;
      memory_array[4411] <= 3'b000;
      memory_array[4412] <= 3'b000;
      memory_array[4413] <= 3'b110;
      memory_array[4414] <= 3'b110;
      memory_array[4415] <= 3'b000;
      memory_array[4416] <= 3'b101;
      memory_array[4417] <= 3'b000;
      memory_array[4418] <= 3'b000;
      memory_array[4419] <= 3'b000;
      memory_array[4420] <= 3'b101;
      memory_array[4421] <= 3'b000;
      memory_array[4422] <= 3'b000;
      memory_array[4423] <= 3'b000;
      memory_array[4424] <= 3'b000;
      memory_array[4425] <= 3'b000;
      memory_array[4426] <= 3'b000;
      memory_array[4427] <= 3'b000;
      memory_array[4428] <= 3'b110;
      memory_array[4429] <= 3'b110;
      memory_array[4430] <= 3'b000;
      memory_array[4431] <= 3'b000;
      memory_array[4432] <= 3'b101;
      memory_array[4433] <= 3'b101;
      memory_array[4434] <= 3'b000;
      memory_array[4435] <= 3'b000;
      memory_array[4436] <= 3'b000;
      memory_array[4437] <= 3'b000;
      memory_array[4438] <= 3'b110;
      memory_array[4439] <= 3'b110;
      memory_array[4440] <= 3'b000;
      memory_array[4441] <= 3'b000;
      memory_array[4442] <= 3'b000;
      memory_array[4443] <= 3'b110;
      memory_array[4444] <= 3'b101;
      memory_array[4445] <= 3'b101;
      memory_array[4446] <= 3'b111;
      memory_array[4447] <= 3'b101;
      memory_array[4448] <= 3'b000;
      memory_array[4449] <= 3'b101;
      memory_array[4450] <= 3'b000;
      memory_array[4451] <= 3'b101;
      memory_array[4452] <= 3'b000;
      memory_array[4453] <= 3'b101;
      memory_array[4454] <= 3'b000;
      memory_array[4455] <= 3'b101;
      memory_array[4456] <= 3'b000;
      memory_array[4457] <= 3'b111;
      memory_array[4458] <= 3'b111;
      memory_array[4459] <= 3'b111;
      memory_array[4460] <= 3'b111;
      memory_array[4461] <= 3'b111;
      memory_array[4462] <= 3'b111;
      memory_array[4463] <= 3'b111;
      memory_array[4464] <= 3'b111;
      memory_array[4465] <= 3'b101;
      memory_array[4466] <= 3'b000;
      memory_array[4467] <= 3'b000;
      memory_array[4468] <= 3'b101;
      memory_array[4469] <= 3'b101;
      memory_array[4470] <= 3'b000;
      memory_array[4471] <= 3'b101;
      memory_array[4472] <= 3'b101;
      memory_array[4473] <= 3'b101;
      memory_array[4474] <= 3'b101;
      memory_array[4475] <= 3'b000;
      memory_array[4476] <= 3'b000;
      memory_array[4477] <= 3'b000;
      memory_array[4478] <= 3'b101;
      memory_array[4479] <= 3'b101;
      memory_array[4480] <= 3'b000;
      memory_array[4481] <= 3'b101;
      memory_array[4482] <= 3'b101;
      memory_array[4483] <= 3'b000;
      memory_array[4484] <= 3'b101;
      memory_array[4485] <= 3'b000;
      memory_array[4486] <= 3'b000;
      memory_array[4487] <= 3'b101;
      memory_array[4488] <= 3'b000;
      memory_array[4489] <= 3'b101;
      memory_array[4490] <= 3'b000;
      memory_array[4491] <= 3'b000;
      memory_array[4492] <= 3'b000;
      memory_array[4493] <= 3'b000;
      memory_array[4494] <= 3'b000;
      memory_array[4495] <= 3'b000;
      memory_array[4496] <= 3'b000;
      memory_array[4497] <= 3'b101;
      memory_array[4498] <= 3'b101;
      memory_array[4499] <= 3'b101;
      memory_array[4500] <= 3'b000;
      memory_array[4501] <= 3'b000;
      memory_array[4502] <= 3'b000;
      memory_array[4503] <= 3'b101;
      memory_array[4504] <= 3'b000;
      memory_array[4505] <= 3'b000;
      memory_array[4506] <= 3'b000;
      memory_array[4507] <= 3'b000;
      memory_array[4508] <= 3'b000;
      memory_array[4509] <= 3'b101;
      memory_array[4510] <= 3'b000;
      memory_array[4511] <= 3'b000;
      memory_array[4512] <= 3'b000;
      memory_array[4513] <= 3'b101;
      memory_array[4514] <= 3'b101;
      memory_array[4515] <= 3'b000;
      memory_array[4516] <= 3'b000;
      memory_array[4517] <= 3'b000;
      memory_array[4518] <= 3'b000;
      memory_array[4519] <= 3'b101;
      memory_array[4520] <= 3'b101;
      memory_array[4521] <= 3'b000;
      memory_array[4522] <= 3'b000;
      memory_array[4523] <= 3'b000;
      memory_array[4524] <= 3'b000;
      memory_array[4525] <= 3'b101;
      memory_array[4526] <= 3'b000;
      memory_array[4527] <= 3'b000;
      memory_array[4528] <= 3'b101;
      memory_array[4529] <= 3'b000;
      memory_array[4530] <= 3'b000;
      memory_array[4531] <= 3'b101;
      memory_array[4532] <= 3'b000;
      memory_array[4533] <= 3'b000;
      memory_array[4534] <= 3'b101;
      memory_array[4535] <= 3'b111;
      memory_array[4536] <= 3'b111;
      memory_array[4537] <= 3'b111;
      memory_array[4538] <= 3'b111;
      memory_array[4539] <= 3'b111;
      memory_array[4540] <= 3'b111;
      memory_array[4541] <= 3'b111;
      memory_array[4542] <= 3'b101;
      memory_array[4543] <= 3'b000;
      memory_array[4544] <= 3'b101;
      memory_array[4545] <= 3'b000;
      memory_array[4546] <= 3'b101;
      memory_array[4547] <= 3'b000;
      memory_array[4548] <= 3'b101;
      memory_array[4549] <= 3'b000;
      memory_array[4550] <= 3'b101;
      memory_array[4551] <= 3'b000;
      memory_array[4552] <= 3'b000;
      memory_array[4553] <= 3'b111;
      memory_array[4554] <= 3'b101;
      memory_array[4555] <= 3'b101;
      memory_array[4556] <= 3'b000;
      memory_array[4557] <= 3'b000;
      memory_array[4558] <= 3'b110;
      memory_array[4559] <= 3'b110;
      memory_array[4560] <= 3'b000;
      memory_array[4561] <= 3'b000;
      memory_array[4562] <= 3'b000;
      memory_array[4563] <= 3'b110;
      memory_array[4564] <= 3'b110;
      memory_array[4565] <= 3'b000;
      memory_array[4566] <= 3'b101;
      memory_array[4567] <= 3'b000;
      memory_array[4568] <= 3'b110;
      memory_array[4569] <= 3'b110;
      memory_array[4570] <= 3'b000;
      memory_array[4571] <= 3'b000;
      memory_array[4572] <= 3'b000;
      memory_array[4573] <= 3'b110;
      memory_array[4574] <= 3'b000;
      memory_array[4575] <= 3'b000;
      memory_array[4576] <= 3'b000;
      memory_array[4577] <= 3'b000;
      memory_array[4578] <= 3'b110;
      memory_array[4579] <= 3'b101;
      memory_array[4580] <= 3'b000;
      memory_array[4581] <= 3'b000;
      memory_array[4582] <= 3'b000;
      memory_array[4583] <= 3'b101;
      memory_array[4584] <= 3'b110;
      memory_array[4585] <= 3'b000;
      memory_array[4586] <= 3'b000;
      memory_array[4587] <= 3'b000;
      memory_array[4588] <= 3'b110;
      memory_array[4589] <= 3'b000;
      memory_array[4590] <= 3'b000;
      memory_array[4591] <= 3'b101;
      memory_array[4592] <= 3'b101;
      memory_array[4593] <= 3'b101;
      memory_array[4594] <= 3'b101;
      memory_array[4595] <= 3'b101;
      memory_array[4596] <= 3'b101;
      memory_array[4597] <= 3'b101;
      memory_array[4598] <= 3'b101;
      memory_array[4599] <= 3'b101;
      memory_array[4600] <= 3'b101;
      memory_array[4601] <= 3'b101;
      memory_array[4602] <= 3'b101;
      memory_array[4603] <= 3'b101;
      memory_array[4604] <= 3'b101;
      memory_array[4605] <= 3'b101;
      memory_array[4606] <= 3'b101;
      memory_array[4607] <= 3'b101;
      memory_array[4608] <= 3'b101;
      memory_array[4609] <= 3'b000;
      memory_array[4610] <= 3'b000;
      memory_array[4611] <= 3'b110;
      memory_array[4612] <= 3'b000;
      memory_array[4613] <= 3'b101;
      memory_array[4614] <= 3'b101;
      memory_array[4615] <= 3'b000;
      memory_array[4616] <= 3'b000;
      memory_array[4617] <= 3'b111;
      memory_array[4618] <= 3'b000;
      memory_array[4619] <= 3'b101;
      memory_array[4620] <= 3'b000;
      memory_array[4621] <= 3'b110;
      memory_array[4622] <= 3'b000;
      memory_array[4623] <= 3'b000;
      memory_array[4624] <= 3'b101;
      memory_array[4625] <= 3'b000;
      memory_array[4626] <= 3'b110;
      memory_array[4627] <= 3'b110;
      memory_array[4628] <= 3'b000;
      memory_array[4629] <= 3'b000;
      memory_array[4630] <= 3'b110;
      memory_array[4631] <= 3'b000;
      memory_array[4632] <= 3'b101;
      memory_array[4633] <= 3'b000;
      memory_array[4634] <= 3'b101;
      memory_array[4635] <= 3'b000;
      memory_array[4636] <= 3'b000;
      memory_array[4637] <= 3'b101;
      memory_array[4638] <= 3'b000;
      memory_array[4639] <= 3'b000;
      memory_array[4640] <= 3'b110;
      memory_array[4641] <= 3'b110;
      memory_array[4642] <= 3'b110;
      memory_array[4643] <= 3'b000;
      memory_array[4644] <= 3'b000;
      memory_array[4645] <= 3'b000;
      memory_array[4646] <= 3'b000;
      memory_array[4647] <= 3'b000;
      memory_array[4648] <= 3'b101;
      memory_array[4649] <= 3'b000;
      memory_array[4650] <= 3'b110;
      memory_array[4651] <= 3'b110;
      memory_array[4652] <= 3'b000;
      memory_array[4653] <= 3'b000;
      memory_array[4654] <= 3'b000;
      memory_array[4655] <= 3'b000;
      memory_array[4656] <= 3'b111;
      memory_array[4657] <= 3'b111;
      memory_array[4658] <= 3'b111;
      memory_array[4659] <= 3'b111;
      memory_array[4660] <= 3'b111;
      memory_array[4661] <= 3'b111;
      memory_array[4662] <= 3'b111;
      memory_array[4663] <= 3'b111;
      memory_array[4664] <= 3'b000;
      memory_array[4665] <= 3'b000;
      memory_array[4666] <= 3'b101;
      memory_array[4667] <= 3'b000;
      memory_array[4668] <= 3'b101;
      memory_array[4669] <= 3'b000;
      memory_array[4670] <= 3'b101;
      memory_array[4671] <= 3'b101;
      memory_array[4672] <= 3'b101;
      memory_array[4673] <= 3'b000;
      memory_array[4674] <= 3'b000;
      memory_array[4675] <= 3'b101;
      memory_array[4676] <= 3'b000;
      memory_array[4677] <= 3'b000;
      memory_array[4678] <= 3'b101;
      memory_array[4679] <= 3'b000;
      memory_array[4680] <= 3'b101;
      memory_array[4681] <= 3'b101;
      memory_array[4682] <= 3'b000;
      memory_array[4683] <= 3'b000;
      memory_array[4684] <= 3'b000;
      memory_array[4685] <= 3'b101;
      memory_array[4686] <= 3'b101;
      memory_array[4687] <= 3'b101;
      memory_array[4688] <= 3'b000;
      memory_array[4689] <= 3'b000;
      memory_array[4690] <= 3'b101;
      memory_array[4691] <= 3'b000;
      memory_array[4692] <= 3'b101;
      memory_array[4693] <= 3'b000;
      memory_array[4694] <= 3'b000;
      memory_array[4695] <= 3'b000;
      memory_array[4696] <= 3'b101;
      memory_array[4697] <= 3'b101;
      memory_array[4698] <= 3'b000;
      memory_array[4699] <= 3'b000;
      memory_array[4700] <= 3'b101;
      memory_array[4701] <= 3'b000;
      memory_array[4702] <= 3'b101;
      memory_array[4703] <= 3'b000;
      memory_array[4704] <= 3'b000;
      memory_array[4705] <= 3'b000;
      memory_array[4706] <= 3'b000;
      memory_array[4707] <= 3'b101;
      memory_array[4708] <= 3'b000;
      memory_array[4709] <= 3'b000;
      memory_array[4710] <= 3'b000;
      memory_array[4711] <= 3'b000;
      memory_array[4712] <= 3'b101;
      memory_array[4713] <= 3'b000;
      memory_array[4714] <= 3'b101;
      memory_array[4715] <= 3'b101;
      memory_array[4716] <= 3'b101;
      memory_array[4717] <= 3'b101;
      memory_array[4718] <= 3'b000;
      memory_array[4719] <= 3'b101;
      memory_array[4720] <= 3'b111;
      memory_array[4721] <= 3'b101;
      memory_array[4722] <= 3'b101;
      memory_array[4723] <= 3'b000;
      memory_array[4724] <= 3'b000;
      memory_array[4725] <= 3'b000;
      memory_array[4726] <= 3'b000;
      memory_array[4727] <= 3'b101;
      memory_array[4728] <= 3'b000;
      memory_array[4729] <= 3'b000;
      memory_array[4730] <= 3'b000;
      memory_array[4731] <= 3'b101;
      memory_array[4732] <= 3'b000;
      memory_array[4733] <= 3'b101;
      memory_array[4734] <= 3'b000;
      memory_array[4735] <= 3'b000;
      memory_array[4736] <= 3'b111;
      memory_array[4737] <= 3'b111;
      memory_array[4738] <= 3'b111;
      memory_array[4739] <= 3'b111;
      memory_array[4740] <= 3'b111;
      memory_array[4741] <= 3'b111;
      memory_array[4742] <= 3'b111;
      memory_array[4743] <= 3'b111;
      memory_array[4744] <= 3'b000;
      memory_array[4745] <= 3'b000;
      memory_array[4746] <= 3'b000;
      memory_array[4747] <= 3'b110;
      memory_array[4748] <= 3'b000;
      memory_array[4749] <= 3'b000;
      memory_array[4750] <= 3'b110;
      memory_array[4751] <= 3'b101;
      memory_array[4752] <= 3'b101;
      memory_array[4753] <= 3'b000;
      memory_array[4754] <= 3'b000;
      memory_array[4755] <= 3'b000;
      memory_array[4756] <= 3'b110;
      memory_array[4757] <= 3'b110;
      memory_array[4758] <= 3'b000;
      memory_array[4759] <= 3'b000;
      memory_array[4760] <= 3'b110;
      memory_array[4761] <= 3'b000;
      memory_array[4762] <= 3'b101;
      memory_array[4763] <= 3'b000;
      memory_array[4764] <= 3'b000;
      memory_array[4765] <= 3'b101;
      memory_array[4766] <= 3'b000;
      memory_array[4767] <= 3'b101;
      memory_array[4768] <= 3'b000;
      memory_array[4769] <= 3'b000;
      memory_array[4770] <= 3'b110;
      memory_array[4771] <= 3'b110;
      memory_array[4772] <= 3'b110;
      memory_array[4773] <= 3'b000;
      memory_array[4774] <= 3'b000;
      memory_array[4775] <= 3'b101;
      memory_array[4776] <= 3'b000;
      memory_array[4777] <= 3'b000;
      memory_array[4778] <= 3'b000;
      memory_array[4779] <= 3'b000;
      memory_array[4780] <= 3'b101;
      memory_array[4781] <= 3'b000;
      memory_array[4782] <= 3'b000;
      memory_array[4783] <= 3'b000;
      memory_array[4784] <= 3'b000;
      memory_array[4785] <= 3'b101;
      memory_array[4786] <= 3'b101;
      memory_array[4787] <= 3'b000;
      memory_array[4788] <= 3'b000;
      memory_array[4789] <= 3'b000;
      memory_array[4790] <= 3'b000;
      memory_array[4791] <= 3'b101;
      memory_array[4792] <= 3'b101;
      memory_array[4793] <= 3'b101;
      memory_array[4794] <= 3'b101;
      memory_array[4795] <= 3'b101;
      memory_array[4796] <= 3'b101;
      memory_array[4797] <= 3'b101;
      memory_array[4798] <= 3'b101;
      memory_array[4799] <= 3'b101;
      memory_array[4800] <= 3'b000;
      memory_array[4801] <= 3'b000;
      memory_array[4802] <= 3'b000;
      memory_array[4803] <= 3'b110;
      memory_array[4804] <= 3'b110;
      memory_array[4805] <= 3'b000;
      memory_array[4806] <= 3'b000;
      memory_array[4807] <= 3'b000;
      memory_array[4808] <= 3'b101;
      memory_array[4809] <= 3'b000;
      memory_array[4810] <= 3'b000;
      memory_array[4811] <= 3'b000;
      memory_array[4812] <= 3'b101;
      memory_array[4813] <= 3'b101;
      memory_array[4814] <= 3'b000;
      memory_array[4815] <= 3'b101;
      memory_array[4816] <= 3'b000;
      memory_array[4817] <= 3'b000;
      memory_array[4818] <= 3'b111;
      memory_array[4819] <= 3'b110;
      memory_array[4820] <= 3'b000;
      memory_array[4821] <= 3'b000;
      memory_array[4822] <= 3'b000;
      memory_array[4823] <= 3'b000;
      memory_array[4824] <= 3'b000;
      memory_array[4825] <= 3'b000;
      memory_array[4826] <= 3'b000;
      memory_array[4827] <= 3'b000;
      memory_array[4828] <= 3'b110;
      memory_array[4829] <= 3'b110;
      memory_array[4830] <= 3'b000;
      memory_array[4831] <= 3'b101;
      memory_array[4832] <= 3'b000;
      memory_array[4833] <= 3'b101;
      memory_array[4834] <= 3'b101;
      memory_array[4835] <= 3'b101;
      memory_array[4836] <= 3'b101;
      memory_array[4837] <= 3'b000;
      memory_array[4838] <= 3'b101;
      memory_array[4839] <= 3'b110;
      memory_array[4840] <= 3'b000;
      memory_array[4841] <= 3'b000;
      memory_array[4842] <= 3'b000;
      memory_array[4843] <= 3'b110;
      memory_array[4844] <= 3'b110;
      memory_array[4845] <= 3'b000;
      memory_array[4846] <= 3'b101;
      memory_array[4847] <= 3'b101;
      memory_array[4848] <= 3'b000;
      memory_array[4849] <= 3'b000;
      memory_array[4850] <= 3'b000;
      memory_array[4851] <= 3'b000;
      memory_array[4852] <= 3'b101;
      memory_array[4853] <= 3'b000;
      memory_array[4854] <= 3'b101;
      memory_array[4855] <= 3'b111;
      memory_array[4856] <= 3'b111;
      memory_array[4857] <= 3'b111;
      memory_array[4858] <= 3'b111;
      memory_array[4859] <= 3'b111;
      memory_array[4860] <= 3'b111;
      memory_array[4861] <= 3'b111;
      memory_array[4862] <= 3'b101;
      memory_array[4863] <= 3'b000;
      memory_array[4864] <= 3'b101;
      memory_array[4865] <= 3'b000;
      memory_array[4866] <= 3'b000;
      memory_array[4867] <= 3'b000;
      memory_array[4868] <= 3'b101;
      memory_array[4869] <= 3'b101;
      memory_array[4870] <= 3'b000;
      memory_array[4871] <= 3'b101;
      memory_array[4872] <= 3'b000;
      memory_array[4873] <= 3'b101;
      memory_array[4874] <= 3'b101;
      memory_array[4875] <= 3'b000;
      memory_array[4876] <= 3'b000;
      memory_array[4877] <= 3'b000;
      memory_array[4878] <= 3'b000;
      memory_array[4879] <= 3'b101;
      memory_array[4880] <= 3'b101;
      memory_array[4881] <= 3'b000;
      memory_array[4882] <= 3'b000;
      memory_array[4883] <= 3'b101;
      memory_array[4884] <= 3'b000;
      memory_array[4885] <= 3'b000;
      memory_array[4886] <= 3'b000;
      memory_array[4887] <= 3'b000;
      memory_array[4888] <= 3'b101;
      memory_array[4889] <= 3'b000;
      memory_array[4890] <= 3'b000;
      memory_array[4891] <= 3'b101;
      memory_array[4892] <= 3'b000;
      memory_array[4893] <= 3'b000;
      memory_array[4894] <= 3'b000;
      memory_array[4895] <= 3'b101;
      memory_array[4896] <= 3'b000;
      memory_array[4897] <= 3'b101;
      memory_array[4898] <= 3'b000;
      memory_array[4899] <= 3'b101;
      memory_array[4900] <= 3'b101;
      memory_array[4901] <= 3'b000;
      memory_array[4902] <= 3'b000;
      memory_array[4903] <= 3'b101;
      memory_array[4904] <= 3'b000;
      memory_array[4905] <= 3'b101;
      memory_array[4906] <= 3'b101;
      memory_array[4907] <= 3'b000;
      memory_array[4908] <= 3'b000;
      memory_array[4909] <= 3'b101;
      memory_array[4910] <= 3'b000;
      memory_array[4911] <= 3'b000;
      memory_array[4912] <= 3'b000;
      memory_array[4913] <= 3'b101;
      memory_array[4914] <= 3'b000;
      memory_array[4915] <= 3'b000;
      memory_array[4916] <= 3'b101;
      memory_array[4917] <= 3'b000;
      memory_array[4918] <= 3'b101;
      memory_array[4919] <= 3'b101;
      memory_array[4920] <= 3'b101;
      memory_array[4921] <= 3'b000;
      memory_array[4922] <= 3'b000;
      memory_array[4923] <= 3'b000;
      memory_array[4924] <= 3'b101;
      memory_array[4925] <= 3'b000;
      memory_array[4926] <= 3'b000;
      memory_array[4927] <= 3'b000;
      memory_array[4928] <= 3'b101;
      memory_array[4929] <= 3'b101;
      memory_array[4930] <= 3'b000;
      memory_array[4931] <= 3'b000;
      memory_array[4932] <= 3'b000;
      memory_array[4933] <= 3'b000;
      memory_array[4934] <= 3'b000;
      memory_array[4935] <= 3'b000;
      memory_array[4936] <= 3'b000;
      memory_array[4937] <= 3'b111;
      memory_array[4938] <= 3'b111;
      memory_array[4939] <= 3'b111;
      memory_array[4940] <= 3'b111;
      memory_array[4941] <= 3'b111;
      memory_array[4942] <= 3'b111;
      memory_array[4943] <= 3'b111;
      memory_array[4944] <= 3'b111;
      memory_array[4945] <= 3'b101;
      memory_array[4946] <= 3'b000;
      memory_array[4947] <= 3'b000;
      memory_array[4948] <= 3'b000;
      memory_array[4949] <= 3'b000;
      memory_array[4950] <= 3'b000;
      memory_array[4951] <= 3'b000;
      memory_array[4952] <= 3'b111;
      memory_array[4953] <= 3'b101;
      memory_array[4954] <= 3'b000;
      memory_array[4955] <= 3'b000;
      memory_array[4956] <= 3'b000;
      memory_array[4957] <= 3'b000;
      memory_array[4958] <= 3'b110;
      memory_array[4959] <= 3'b110;
      memory_array[4960] <= 3'b000;
      memory_array[4961] <= 3'b101;
      memory_array[4962] <= 3'b000;
      memory_array[4963] <= 3'b101;
      memory_array[4964] <= 3'b101;
      memory_array[4965] <= 3'b101;
      memory_array[4966] <= 3'b101;
      memory_array[4967] <= 3'b101;
      memory_array[4968] <= 3'b101;
      memory_array[4969] <= 3'b110;
      memory_array[4970] <= 3'b000;
      memory_array[4971] <= 3'b000;
      memory_array[4972] <= 3'b000;
      memory_array[4973] <= 3'b110;
      memory_array[4974] <= 3'b110;
      memory_array[4975] <= 3'b000;
      memory_array[4976] <= 3'b000;
      memory_array[4977] <= 3'b000;
      memory_array[4978] <= 3'b110;
      memory_array[4979] <= 3'b000;
      memory_array[4980] <= 3'b111;
      memory_array[4981] <= 3'b111;
      memory_array[4982] <= 3'b000;
      memory_array[4983] <= 3'b000;
      memory_array[4984] <= 3'b101;
      memory_array[4985] <= 3'b000;
      memory_array[4986] <= 3'b101;
      memory_array[4987] <= 3'b000;
      memory_array[4988] <= 3'b110;
      memory_array[4989] <= 3'b000;
      memory_array[4990] <= 3'b000;
      memory_array[4991] <= 3'b101;
      memory_array[4992] <= 3'b000;
      memory_array[4993] <= 3'b110;
      memory_array[4994] <= 3'b110;
      memory_array[4995] <= 3'b000;
      memory_array[4996] <= 3'b000;
      memory_array[4997] <= 3'b000;
      memory_array[4998] <= 3'b110;
      memory_array[4999] <= 3'b110;
      memory_array[5000] <= 3'b101;
      memory_array[5001] <= 3'b110;
      memory_array[5002] <= 3'b110;
      memory_array[5003] <= 3'b000;
      memory_array[5004] <= 3'b000;
      memory_array[5005] <= 3'b110;
      memory_array[5006] <= 3'b110;
      memory_array[5007] <= 3'b101;
      memory_array[5008] <= 3'b101;
      memory_array[5009] <= 3'b000;
      memory_array[5010] <= 3'b000;
      memory_array[5011] <= 3'b110;
      memory_array[5012] <= 3'b101;
      memory_array[5013] <= 3'b000;
      memory_array[5014] <= 3'b000;
      memory_array[5015] <= 3'b101;
      memory_array[5016] <= 3'b000;
      memory_array[5017] <= 3'b111;
      memory_array[5018] <= 3'b000;
      memory_array[5019] <= 3'b101;
      memory_array[5020] <= 3'b000;
      memory_array[5021] <= 3'b110;
      memory_array[5022] <= 3'b101;
      memory_array[5023] <= 3'b101;
      memory_array[5024] <= 3'b000;
      memory_array[5025] <= 3'b110;
      memory_array[5026] <= 3'b110;
      memory_array[5027] <= 3'b110;
      memory_array[5028] <= 3'b000;
      memory_array[5029] <= 3'b000;
      memory_array[5030] <= 3'b110;
      memory_array[5031] <= 3'b000;
      memory_array[5032] <= 3'b101;
      memory_array[5033] <= 3'b000;
      memory_array[5034] <= 3'b101;
      memory_array[5035] <= 3'b000;
      memory_array[5036] <= 3'b110;
      memory_array[5037] <= 3'b000;
      memory_array[5038] <= 3'b101;
      memory_array[5039] <= 3'b000;
      memory_array[5040] <= 3'b110;
      memory_array[5041] <= 3'b110;
      memory_array[5042] <= 3'b110;
      memory_array[5043] <= 3'b000;
      memory_array[5044] <= 3'b000;
      memory_array[5045] <= 3'b000;
      memory_array[5046] <= 3'b000;
      memory_array[5047] <= 3'b000;
      memory_array[5048] <= 3'b101;
      memory_array[5049] <= 3'b000;
      memory_array[5050] <= 3'b000;
      memory_array[5051] <= 3'b000;
      memory_array[5052] <= 3'b000;
      memory_array[5053] <= 3'b101;
      memory_array[5054] <= 3'b111;
      memory_array[5055] <= 3'b111;
      memory_array[5056] <= 3'b111;
      memory_array[5057] <= 3'b111;
      memory_array[5058] <= 3'b111;
      memory_array[5059] <= 3'b111;
      memory_array[5060] <= 3'b111;
      memory_array[5061] <= 3'b000;
      memory_array[5062] <= 3'b000;
      memory_array[5063] <= 3'b000;
      memory_array[5064] <= 3'b101;
      memory_array[5065] <= 3'b101;
      memory_array[5066] <= 3'b101;
      memory_array[5067] <= 3'b000;
      memory_array[5068] <= 3'b000;
      memory_array[5069] <= 3'b000;
      memory_array[5070] <= 3'b101;
      memory_array[5071] <= 3'b101;
      memory_array[5072] <= 3'b000;
      memory_array[5073] <= 3'b000;
      memory_array[5074] <= 3'b000;
      memory_array[5075] <= 3'b101;
      memory_array[5076] <= 3'b000;
      memory_array[5077] <= 3'b101;
      memory_array[5078] <= 3'b000;
      memory_array[5079] <= 3'b000;
      memory_array[5080] <= 3'b000;
      memory_array[5081] <= 3'b101;
      memory_array[5082] <= 3'b101;
      memory_array[5083] <= 3'b101;
      memory_array[5084] <= 3'b000;
      memory_array[5085] <= 3'b000;
      memory_array[5086] <= 3'b101;
      memory_array[5087] <= 3'b101;
      memory_array[5088] <= 3'b000;
      memory_array[5089] <= 3'b000;
      memory_array[5090] <= 3'b101;
      memory_array[5091] <= 3'b000;
      memory_array[5092] <= 3'b101;
      memory_array[5093] <= 3'b000;
      memory_array[5094] <= 3'b101;
      memory_array[5095] <= 3'b000;
      memory_array[5096] <= 3'b000;
      memory_array[5097] <= 3'b000;
      memory_array[5098] <= 3'b000;
      memory_array[5099] <= 3'b000;
      memory_array[5100] <= 3'b000;
      memory_array[5101] <= 3'b000;
      memory_array[5102] <= 3'b000;
      memory_array[5103] <= 3'b000;
      memory_array[5104] <= 3'b000;
      memory_array[5105] <= 3'b101;
      memory_array[5106] <= 3'b000;
      memory_array[5107] <= 3'b101;
      memory_array[5108] <= 3'b101;
      memory_array[5109] <= 3'b000;
      memory_array[5110] <= 3'b101;
      memory_array[5111] <= 3'b101;
      memory_array[5112] <= 3'b101;
      memory_array[5113] <= 3'b000;
      memory_array[5114] <= 3'b000;
      memory_array[5115] <= 3'b000;
      memory_array[5116] <= 3'b101;
      memory_array[5117] <= 3'b101;
      memory_array[5118] <= 3'b101;
      memory_array[5119] <= 3'b000;
      memory_array[5120] <= 3'b000;
      memory_array[5121] <= 3'b101;
      memory_array[5122] <= 3'b101;
      memory_array[5123] <= 3'b101;
      memory_array[5124] <= 3'b000;
      memory_array[5125] <= 3'b000;
      memory_array[5126] <= 3'b101;
      memory_array[5127] <= 3'b000;
      memory_array[5128] <= 3'b000;
      memory_array[5129] <= 3'b000;
      memory_array[5130] <= 3'b101;
      memory_array[5131] <= 3'b000;
      memory_array[5132] <= 3'b101;
      memory_array[5133] <= 3'b000;
      memory_array[5134] <= 3'b000;
      memory_array[5135] <= 3'b101;
      memory_array[5136] <= 3'b101;
      memory_array[5137] <= 3'b000;
      memory_array[5138] <= 3'b000;
      memory_array[5139] <= 3'b111;
      memory_array[5140] <= 3'b111;
      memory_array[5141] <= 3'b111;
      memory_array[5142] <= 3'b111;
      memory_array[5143] <= 3'b111;
      memory_array[5144] <= 3'b111;
      memory_array[5145] <= 3'b111;
      memory_array[5146] <= 3'b101;
      memory_array[5147] <= 3'b000;
      memory_array[5148] <= 3'b000;
      memory_array[5149] <= 3'b000;
      memory_array[5150] <= 3'b000;
      memory_array[5151] <= 3'b101;
      memory_array[5152] <= 3'b101;
      memory_array[5153] <= 3'b000;
      memory_array[5154] <= 3'b000;
      memory_array[5155] <= 3'b110;
      memory_array[5156] <= 3'b110;
      memory_array[5157] <= 3'b110;
      memory_array[5158] <= 3'b000;
      memory_array[5159] <= 3'b000;
      memory_array[5160] <= 3'b110;
      memory_array[5161] <= 3'b101;
      memory_array[5162] <= 3'b110;
      memory_array[5163] <= 3'b000;
      memory_array[5164] <= 3'b000;
      memory_array[5165] <= 3'b101;
      memory_array[5166] <= 3'b000;
      memory_array[5167] <= 3'b101;
      memory_array[5168] <= 3'b000;
      memory_array[5169] <= 3'b000;
      memory_array[5170] <= 3'b110;
      memory_array[5171] <= 3'b110;
      memory_array[5172] <= 3'b110;
      memory_array[5173] <= 3'b000;
      memory_array[5174] <= 3'b000;
      memory_array[5175] <= 3'b110;
      memory_array[5176] <= 3'b101;
      memory_array[5177] <= 3'b000;
      memory_array[5178] <= 3'b000;
      memory_array[5179] <= 3'b000;
      memory_array[5180] <= 3'b101;
      memory_array[5181] <= 3'b000;
      memory_array[5182] <= 3'b000;
      memory_array[5183] <= 3'b000;
      memory_array[5184] <= 3'b101;
      memory_array[5185] <= 3'b000;
      memory_array[5186] <= 3'b000;
      memory_array[5187] <= 3'b000;
      memory_array[5188] <= 3'b000;
      memory_array[5189] <= 3'b000;
      memory_array[5190] <= 3'b000;
      memory_array[5191] <= 3'b101;
      memory_array[5192] <= 3'b110;
      memory_array[5193] <= 3'b000;
      memory_array[5194] <= 3'b000;
      memory_array[5195] <= 3'b110;
      memory_array[5196] <= 3'b110;
      memory_array[5197] <= 3'b110;
      memory_array[5198] <= 3'b000;
      memory_array[5199] <= 3'b101;
      memory_array[5200] <= 3'b101;
      memory_array[5201] <= 3'b101;
      memory_array[5202] <= 3'b110;
      memory_array[5203] <= 3'b101;
      memory_array[5204] <= 3'b101;
      memory_array[5205] <= 3'b110;
      memory_array[5206] <= 3'b101;
      memory_array[5207] <= 3'b101;
      memory_array[5208] <= 3'b101;
      memory_array[5209] <= 3'b000;
      memory_array[5210] <= 3'b000;
      memory_array[5211] <= 3'b110;
      memory_array[5212] <= 3'b101;
      memory_array[5213] <= 3'b000;
      memory_array[5214] <= 3'b000;
      memory_array[5215] <= 3'b110;
      memory_array[5216] <= 3'b110;
      memory_array[5217] <= 3'b000;
      memory_array[5218] <= 3'b000;
      memory_array[5219] <= 3'b000;
      memory_array[5220] <= 3'b110;
      memory_array[5221] <= 3'b110;
      memory_array[5222] <= 3'b110;
      memory_array[5223] <= 3'b000;
      memory_array[5224] <= 3'b000;
      memory_array[5225] <= 3'b101;
      memory_array[5226] <= 3'b101;
      memory_array[5227] <= 3'b110;
      memory_array[5228] <= 3'b000;
      memory_array[5229] <= 3'b000;
      memory_array[5230] <= 3'b110;
      memory_array[5231] <= 3'b110;
      memory_array[5232] <= 3'b000;
      memory_array[5233] <= 3'b101;
      memory_array[5234] <= 3'b000;
      memory_array[5235] <= 3'b110;
      memory_array[5236] <= 3'b110;
      memory_array[5237] <= 3'b110;
      memory_array[5238] <= 3'b000;
      memory_array[5239] <= 3'b000;
      memory_array[5240] <= 3'b110;
      memory_array[5241] <= 3'b110;
      memory_array[5242] <= 3'b110;
      memory_array[5243] <= 3'b000;
      memory_array[5244] <= 3'b000;
      memory_array[5245] <= 3'b000;
      memory_array[5246] <= 3'b000;
      memory_array[5247] <= 3'b000;
      memory_array[5248] <= 3'b101;
      memory_array[5249] <= 3'b000;
      memory_array[5250] <= 3'b000;
      memory_array[5251] <= 3'b101;
      memory_array[5252] <= 3'b111;
      memory_array[5253] <= 3'b111;
      memory_array[5254] <= 3'b111;
      memory_array[5255] <= 3'b111;
      memory_array[5256] <= 3'b111;
      memory_array[5257] <= 3'b111;
      memory_array[5258] <= 3'b101;
      memory_array[5259] <= 3'b000;
      memory_array[5260] <= 3'b101;
      memory_array[5261] <= 3'b000;
      memory_array[5262] <= 3'b101;
      memory_array[5263] <= 3'b000;
      memory_array[5264] <= 3'b000;
      memory_array[5265] <= 3'b101;
      memory_array[5266] <= 3'b101;
      memory_array[5267] <= 3'b101;
      memory_array[5268] <= 3'b000;
      memory_array[5269] <= 3'b000;
      memory_array[5270] <= 3'b101;
      memory_array[5271] <= 3'b101;
      memory_array[5272] <= 3'b101;
      memory_array[5273] <= 3'b000;
      memory_array[5274] <= 3'b000;
      memory_array[5275] <= 3'b000;
      memory_array[5276] <= 3'b101;
      memory_array[5277] <= 3'b000;
      memory_array[5278] <= 3'b000;
      memory_array[5279] <= 3'b101;
      memory_array[5280] <= 3'b101;
      memory_array[5281] <= 3'b101;
      memory_array[5282] <= 3'b000;
      memory_array[5283] <= 3'b000;
      memory_array[5284] <= 3'b000;
      memory_array[5285] <= 3'b101;
      memory_array[5286] <= 3'b101;
      memory_array[5287] <= 3'b101;
      memory_array[5288] <= 3'b000;
      memory_array[5289] <= 3'b101;
      memory_array[5290] <= 3'b101;
      memory_array[5291] <= 3'b101;
      memory_array[5292] <= 3'b000;
      memory_array[5293] <= 3'b101;
      memory_array[5294] <= 3'b000;
      memory_array[5295] <= 3'b000;
      memory_array[5296] <= 3'b101;
      memory_array[5297] <= 3'b101;
      memory_array[5298] <= 3'b000;
      memory_array[5299] <= 3'b101;
      memory_array[5300] <= 3'b101;
      memory_array[5301] <= 3'b000;
      memory_array[5302] <= 3'b000;
      memory_array[5303] <= 3'b000;
      memory_array[5304] <= 3'b101;
      memory_array[5305] <= 3'b101;
      memory_array[5306] <= 3'b000;
      memory_array[5307] <= 3'b101;
      memory_array[5308] <= 3'b101;
      memory_array[5309] <= 3'b000;
      memory_array[5310] <= 3'b000;
      memory_array[5311] <= 3'b101;
      memory_array[5312] <= 3'b101;
      memory_array[5313] <= 3'b000;
      memory_array[5314] <= 3'b000;
      memory_array[5315] <= 3'b101;
      memory_array[5316] <= 3'b000;
      memory_array[5317] <= 3'b101;
      memory_array[5318] <= 3'b000;
      memory_array[5319] <= 3'b101;
      memory_array[5320] <= 3'b101;
      memory_array[5321] <= 3'b000;
      memory_array[5322] <= 3'b111;
      memory_array[5323] <= 3'b111;
      memory_array[5324] <= 3'b000;
      memory_array[5325] <= 3'b101;
      memory_array[5326] <= 3'b101;
      memory_array[5327] <= 3'b101;
      memory_array[5328] <= 3'b101;
      memory_array[5329] <= 3'b101;
      memory_array[5330] <= 3'b000;
      memory_array[5331] <= 3'b000;
      memory_array[5332] <= 3'b000;
      memory_array[5333] <= 3'b000;
      memory_array[5334] <= 3'b101;
      memory_array[5335] <= 3'b000;
      memory_array[5336] <= 3'b000;
      memory_array[5337] <= 3'b101;
      memory_array[5338] <= 3'b000;
      memory_array[5339] <= 3'b000;
      memory_array[5340] <= 3'b000;
      memory_array[5341] <= 3'b101;
      memory_array[5342] <= 3'b111;
      memory_array[5343] <= 3'b111;
      memory_array[5344] <= 3'b111;
      memory_array[5345] <= 3'b111;
      memory_array[5346] <= 3'b111;
      memory_array[5347] <= 3'b111;
      memory_array[5348] <= 3'b101;
      memory_array[5349] <= 3'b000;
      memory_array[5350] <= 3'b110;
      memory_array[5351] <= 3'b101;
      memory_array[5352] <= 3'b000;
      memory_array[5353] <= 3'b000;
      memory_array[5354] <= 3'b000;
      memory_array[5355] <= 3'b000;
      memory_array[5356] <= 3'b110;
      memory_array[5357] <= 3'b110;
      memory_array[5358] <= 3'b000;
      memory_array[5359] <= 3'b000;
      memory_array[5360] <= 3'b000;
      memory_array[5361] <= 3'b000;
      memory_array[5362] <= 3'b110;
      memory_array[5363] <= 3'b000;
      memory_array[5364] <= 3'b000;
      memory_array[5365] <= 3'b110;
      memory_array[5366] <= 3'b101;
      memory_array[5367] <= 3'b000;
      memory_array[5368] <= 3'b000;
      memory_array[5369] <= 3'b000;
      memory_array[5370] <= 3'b110;
      memory_array[5371] <= 3'b110;
      memory_array[5372] <= 3'b000;
      memory_array[5373] <= 3'b101;
      memory_array[5374] <= 3'b101;
      memory_array[5375] <= 3'b000;
      memory_array[5376] <= 3'b110;
      memory_array[5377] <= 3'b000;
      memory_array[5378] <= 3'b000;
      memory_array[5379] <= 3'b000;
      memory_array[5380] <= 3'b000;
      memory_array[5381] <= 3'b000;
      memory_array[5382] <= 3'b000;
      memory_array[5383] <= 3'b000;
      memory_array[5384] <= 3'b000;
      memory_array[5385] <= 3'b110;
      memory_array[5386] <= 3'b000;
      memory_array[5387] <= 3'b000;
      memory_array[5388] <= 3'b000;
      memory_array[5389] <= 3'b000;
      memory_array[5390] <= 3'b000;
      memory_array[5391] <= 3'b101;
      memory_array[5392] <= 3'b101;
      memory_array[5393] <= 3'b101;
      memory_array[5394] <= 3'b000;
      memory_array[5395] <= 3'b101;
      memory_array[5396] <= 3'b101;
      memory_array[5397] <= 3'b110;
      memory_array[5398] <= 3'b101;
      memory_array[5399] <= 3'b101;
      memory_array[5400] <= 3'b101;
      memory_array[5401] <= 3'b101;
      memory_array[5402] <= 3'b101;
      memory_array[5403] <= 3'b111;
      memory_array[5404] <= 3'b111;
      memory_array[5405] <= 3'b101;
      memory_array[5406] <= 3'b101;
      memory_array[5407] <= 3'b101;
      memory_array[5408] <= 3'b101;
      memory_array[5409] <= 3'b000;
      memory_array[5410] <= 3'b000;
      memory_array[5411] <= 3'b000;
      memory_array[5412] <= 3'b101;
      memory_array[5413] <= 3'b000;
      memory_array[5414] <= 3'b110;
      memory_array[5415] <= 3'b000;
      memory_array[5416] <= 3'b000;
      memory_array[5417] <= 3'b000;
      memory_array[5418] <= 3'b101;
      memory_array[5419] <= 3'b110;
      memory_array[5420] <= 3'b000;
      memory_array[5421] <= 3'b000;
      memory_array[5422] <= 3'b000;
      memory_array[5423] <= 3'b110;
      memory_array[5424] <= 3'b000;
      memory_array[5425] <= 3'b000;
      memory_array[5426] <= 3'b000;
      memory_array[5427] <= 3'b000;
      memory_array[5428] <= 3'b110;
      memory_array[5429] <= 3'b110;
      memory_array[5430] <= 3'b000;
      memory_array[5431] <= 3'b000;
      memory_array[5432] <= 3'b000;
      memory_array[5433] <= 3'b110;
      memory_array[5434] <= 3'b110;
      memory_array[5435] <= 3'b000;
      memory_array[5436] <= 3'b101;
      memory_array[5437] <= 3'b000;
      memory_array[5438] <= 3'b000;
      memory_array[5439] <= 3'b000;
      memory_array[5440] <= 3'b000;
      memory_array[5441] <= 3'b000;
      memory_array[5442] <= 3'b000;
      memory_array[5443] <= 3'b110;
      memory_array[5444] <= 3'b110;
      memory_array[5445] <= 3'b000;
      memory_array[5446] <= 3'b000;
      memory_array[5447] <= 3'b000;
      memory_array[5448] <= 3'b101;
      memory_array[5449] <= 3'b000;
      memory_array[5450] <= 3'b101;
      memory_array[5451] <= 3'b111;
      memory_array[5452] <= 3'b111;
      memory_array[5453] <= 3'b111;
      memory_array[5454] <= 3'b111;
      memory_array[5455] <= 3'b111;
      memory_array[5456] <= 3'b111;
      memory_array[5457] <= 3'b000;
      memory_array[5458] <= 3'b000;
      memory_array[5459] <= 3'b101;
      memory_array[5460] <= 3'b000;
      memory_array[5461] <= 3'b101;
      memory_array[5462] <= 3'b000;
      memory_array[5463] <= 3'b000;
      memory_array[5464] <= 3'b101;
      memory_array[5465] <= 3'b000;
      memory_array[5466] <= 3'b101;
      memory_array[5467] <= 3'b000;
      memory_array[5468] <= 3'b000;
      memory_array[5469] <= 3'b000;
      memory_array[5470] <= 3'b000;
      memory_array[5471] <= 3'b000;
      memory_array[5472] <= 3'b000;
      memory_array[5473] <= 3'b000;
      memory_array[5474] <= 3'b101;
      memory_array[5475] <= 3'b000;
      memory_array[5476] <= 3'b000;
      memory_array[5477] <= 3'b000;
      memory_array[5478] <= 3'b000;
      memory_array[5479] <= 3'b101;
      memory_array[5480] <= 3'b101;
      memory_array[5481] <= 3'b101;
      memory_array[5482] <= 3'b000;
      memory_array[5483] <= 3'b101;
      memory_array[5484] <= 3'b000;
      memory_array[5485] <= 3'b000;
      memory_array[5486] <= 3'b101;
      memory_array[5487] <= 3'b000;
      memory_array[5488] <= 3'b101;
      memory_array[5489] <= 3'b101;
      memory_array[5490] <= 3'b000;
      memory_array[5491] <= 3'b000;
      memory_array[5492] <= 3'b000;
      memory_array[5493] <= 3'b101;
      memory_array[5494] <= 3'b101;
      memory_array[5495] <= 3'b000;
      memory_array[5496] <= 3'b000;
      memory_array[5497] <= 3'b000;
      memory_array[5498] <= 3'b000;
      memory_array[5499] <= 3'b000;
      memory_array[5500] <= 3'b000;
      memory_array[5501] <= 3'b000;
      memory_array[5502] <= 3'b000;
      memory_array[5503] <= 3'b101;
      memory_array[5504] <= 3'b101;
      memory_array[5505] <= 3'b000;
      memory_array[5506] <= 3'b101;
      memory_array[5507] <= 3'b000;
      memory_array[5508] <= 3'b101;
      memory_array[5509] <= 3'b101;
      memory_array[5510] <= 3'b000;
      memory_array[5511] <= 3'b101;
      memory_array[5512] <= 3'b000;
      memory_array[5513] <= 3'b101;
      memory_array[5514] <= 3'b000;
      memory_array[5515] <= 3'b000;
      memory_array[5516] <= 3'b101;
      memory_array[5517] <= 3'b000;
      memory_array[5518] <= 3'b101;
      memory_array[5519] <= 3'b101;
      memory_array[5520] <= 3'b101;
      memory_array[5521] <= 3'b101;
      memory_array[5522] <= 3'b111;
      memory_array[5523] <= 3'b111;
      memory_array[5524] <= 3'b111;
      memory_array[5525] <= 3'b101;
      memory_array[5526] <= 3'b000;
      memory_array[5527] <= 3'b101;
      memory_array[5528] <= 3'b000;
      memory_array[5529] <= 3'b101;
      memory_array[5530] <= 3'b000;
      memory_array[5531] <= 3'b000;
      memory_array[5532] <= 3'b101;
      memory_array[5533] <= 3'b111;
      memory_array[5534] <= 3'b101;
      memory_array[5535] <= 3'b101;
      memory_array[5536] <= 3'b000;
      memory_array[5537] <= 3'b000;
      memory_array[5538] <= 3'b101;
      memory_array[5539] <= 3'b000;
      memory_array[5540] <= 3'b101;
      memory_array[5541] <= 3'b000;
      memory_array[5542] <= 3'b101;
      memory_array[5543] <= 3'b111;
      memory_array[5544] <= 3'b111;
      memory_array[5545] <= 3'b111;
      memory_array[5546] <= 3'b111;
      memory_array[5547] <= 3'b111;
      memory_array[5548] <= 3'b111;
      memory_array[5549] <= 3'b101;
      memory_array[5550] <= 3'b000;
      memory_array[5551] <= 3'b101;
      memory_array[5552] <= 3'b000;
      memory_array[5553] <= 3'b000;
      memory_array[5554] <= 3'b000;
      memory_array[5555] <= 3'b000;
      memory_array[5556] <= 3'b000;
      memory_array[5557] <= 3'b000;
      memory_array[5558] <= 3'b110;
      memory_array[5559] <= 3'b110;
      memory_array[5560] <= 3'b000;
      memory_array[5561] <= 3'b000;
      memory_array[5562] <= 3'b101;
      memory_array[5563] <= 3'b101;
      memory_array[5564] <= 3'b000;
      memory_array[5565] <= 3'b000;
      memory_array[5566] <= 3'b000;
      memory_array[5567] <= 3'b000;
      memory_array[5568] <= 3'b110;
      memory_array[5569] <= 3'b110;
      memory_array[5570] <= 3'b000;
      memory_array[5571] <= 3'b000;
      memory_array[5572] <= 3'b000;
      memory_array[5573] <= 3'b000;
      memory_array[5574] <= 3'b000;
      memory_array[5575] <= 3'b000;
      memory_array[5576] <= 3'b000;
      memory_array[5577] <= 3'b000;
      memory_array[5578] <= 3'b110;
      memory_array[5579] <= 3'b110;
      memory_array[5580] <= 3'b000;
      memory_array[5581] <= 3'b101;
      memory_array[5582] <= 3'b000;
      memory_array[5583] <= 3'b110;
      memory_array[5584] <= 3'b110;
      memory_array[5585] <= 3'b000;
      memory_array[5586] <= 3'b000;
      memory_array[5587] <= 3'b000;
      memory_array[5588] <= 3'b110;
      memory_array[5589] <= 3'b000;
      memory_array[5590] <= 3'b000;
      memory_array[5591] <= 3'b101;
      memory_array[5592] <= 3'b101;
      memory_array[5593] <= 3'b101;
      memory_array[5594] <= 3'b101;
      memory_array[5595] <= 3'b111;
      memory_array[5596] <= 3'b111;
      memory_array[5597] <= 3'b101;
      memory_array[5598] <= 3'b101;
      memory_array[5599] <= 3'b101;
      memory_array[5600] <= 3'b101;
      memory_array[5601] <= 3'b101;
      memory_array[5602] <= 3'b101;
      memory_array[5603] <= 3'b101;
      memory_array[5604] <= 3'b101;
      memory_array[5605] <= 3'b101;
      memory_array[5606] <= 3'b101;
      memory_array[5607] <= 3'b101;
      memory_array[5608] <= 3'b101;
      memory_array[5609] <= 3'b000;
      memory_array[5610] <= 3'b000;
      memory_array[5611] <= 3'b110;
      memory_array[5612] <= 3'b101;
      memory_array[5613] <= 3'b000;
      memory_array[5614] <= 3'b000;
      memory_array[5615] <= 3'b000;
      memory_array[5616] <= 3'b101;
      memory_array[5617] <= 3'b000;
      memory_array[5618] <= 3'b000;
      memory_array[5619] <= 3'b000;
      memory_array[5620] <= 3'b110;
      memory_array[5621] <= 3'b110;
      memory_array[5622] <= 3'b110;
      memory_array[5623] <= 3'b000;
      memory_array[5624] <= 3'b000;
      memory_array[5625] <= 3'b000;
      memory_array[5626] <= 3'b000;
      memory_array[5627] <= 3'b111;
      memory_array[5628] <= 3'b000;
      memory_array[5629] <= 3'b000;
      memory_array[5630] <= 3'b110;
      memory_array[5631] <= 3'b110;
      memory_array[5632] <= 3'b000;
      memory_array[5633] <= 3'b000;
      memory_array[5634] <= 3'b000;
      memory_array[5635] <= 3'b101;
      memory_array[5636] <= 3'b000;
      memory_array[5637] <= 3'b101;
      memory_array[5638] <= 3'b000;
      memory_array[5639] <= 3'b000;
      memory_array[5640] <= 3'b110;
      memory_array[5641] <= 3'b110;
      memory_array[5642] <= 3'b110;
      memory_array[5643] <= 3'b000;
      memory_array[5644] <= 3'b000;
      memory_array[5645] <= 3'b000;
      memory_array[5646] <= 3'b110;
      memory_array[5647] <= 3'b000;
      memory_array[5648] <= 3'b000;
      memory_array[5649] <= 3'b101;
      memory_array[5650] <= 3'b111;
      memory_array[5651] <= 3'b111;
      memory_array[5652] <= 3'b111;
      memory_array[5653] <= 3'b111;
      memory_array[5654] <= 3'b111;
      memory_array[5655] <= 3'b111;
      memory_array[5656] <= 3'b000;
      memory_array[5657] <= 3'b101;
      memory_array[5658] <= 3'b000;
      memory_array[5659] <= 3'b101;
      memory_array[5660] <= 3'b101;
      memory_array[5661] <= 3'b101;
      memory_array[5662] <= 3'b101;
      memory_array[5663] <= 3'b000;
      memory_array[5664] <= 3'b101;
      memory_array[5665] <= 3'b000;
      memory_array[5666] <= 3'b101;
      memory_array[5667] <= 3'b101;
      memory_array[5668] <= 3'b101;
      memory_array[5669] <= 3'b000;
      memory_array[5670] <= 3'b101;
      memory_array[5671] <= 3'b000;
      memory_array[5672] <= 3'b101;
      memory_array[5673] <= 3'b101;
      memory_array[5674] <= 3'b101;
      memory_array[5675] <= 3'b000;
      memory_array[5676] <= 3'b000;
      memory_array[5677] <= 3'b101;
      memory_array[5678] <= 3'b000;
      memory_array[5679] <= 3'b000;
      memory_array[5680] <= 3'b000;
      memory_array[5681] <= 3'b101;
      memory_array[5682] <= 3'b101;
      memory_array[5683] <= 3'b000;
      memory_array[5684] <= 3'b000;
      memory_array[5685] <= 3'b000;
      memory_array[5686] <= 3'b101;
      memory_array[5687] <= 3'b111;
      memory_array[5688] <= 3'b000;
      memory_array[5689] <= 3'b101;
      memory_array[5690] <= 3'b000;
      memory_array[5691] <= 3'b000;
      memory_array[5692] <= 3'b101;
      memory_array[5693] <= 3'b101;
      memory_array[5694] <= 3'b000;
      memory_array[5695] <= 3'b000;
      memory_array[5696] <= 3'b101;
      memory_array[5697] <= 3'b101;
      memory_array[5698] <= 3'b101;
      memory_array[5699] <= 3'b000;
      memory_array[5700] <= 3'b101;
      memory_array[5701] <= 3'b000;
      memory_array[5702] <= 3'b000;
      memory_array[5703] <= 3'b000;
      memory_array[5704] <= 3'b101;
      memory_array[5705] <= 3'b101;
      memory_array[5706] <= 3'b000;
      memory_array[5707] <= 3'b101;
      memory_array[5708] <= 3'b000;
      memory_array[5709] <= 3'b000;
      memory_array[5710] <= 3'b101;
      memory_array[5711] <= 3'b101;
      memory_array[5712] <= 3'b000;
      memory_array[5713] <= 3'b101;
      memory_array[5714] <= 3'b000;
      memory_array[5715] <= 3'b000;
      memory_array[5716] <= 3'b101;
      memory_array[5717] <= 3'b101;
      memory_array[5718] <= 3'b101;
      memory_array[5719] <= 3'b000;
      memory_array[5720] <= 3'b101;
      memory_array[5721] <= 3'b000;
      memory_array[5722] <= 3'b111;
      memory_array[5723] <= 3'b111;
      memory_array[5724] <= 3'b000;
      memory_array[5725] <= 3'b101;
      memory_array[5726] <= 3'b101;
      memory_array[5727] <= 3'b000;
      memory_array[5728] <= 3'b000;
      memory_array[5729] <= 3'b101;
      memory_array[5730] <= 3'b000;
      memory_array[5731] <= 3'b101;
      memory_array[5732] <= 3'b111;
      memory_array[5733] <= 3'b111;
      memory_array[5734] <= 3'b000;
      memory_array[5735] <= 3'b101;
      memory_array[5736] <= 3'b000;
      memory_array[5737] <= 3'b101;
      memory_array[5738] <= 3'b000;
      memory_array[5739] <= 3'b101;
      memory_array[5740] <= 3'b101;
      memory_array[5741] <= 3'b000;
      memory_array[5742] <= 3'b000;
      memory_array[5743] <= 3'b000;
      memory_array[5744] <= 3'b111;
      memory_array[5745] <= 3'b111;
      memory_array[5746] <= 3'b111;
      memory_array[5747] <= 3'b111;
      memory_array[5748] <= 3'b111;
      memory_array[5749] <= 3'b111;
      memory_array[5750] <= 3'b101;
      memory_array[5751] <= 3'b000;
      memory_array[5752] <= 3'b110;
      memory_array[5753] <= 3'b000;
      memory_array[5754] <= 3'b000;
      memory_array[5755] <= 3'b110;
      memory_array[5756] <= 3'b110;
      memory_array[5757] <= 3'b110;
      memory_array[5758] <= 3'b000;
      memory_array[5759] <= 3'b000;
      memory_array[5760] <= 3'b000;
      memory_array[5761] <= 3'b000;
      memory_array[5762] <= 3'b000;
      memory_array[5763] <= 3'b000;
      memory_array[5764] <= 3'b101;
      memory_array[5765] <= 3'b000;
      memory_array[5766] <= 3'b000;
      memory_array[5767] <= 3'b000;
      memory_array[5768] <= 3'b000;
      memory_array[5769] <= 3'b000;
      memory_array[5770] <= 3'b110;
      memory_array[5771] <= 3'b000;
      memory_array[5772] <= 3'b101;
      memory_array[5773] <= 3'b000;
      memory_array[5774] <= 3'b000;
      memory_array[5775] <= 3'b101;
      memory_array[5776] <= 3'b000;
      memory_array[5777] <= 3'b110;
      memory_array[5778] <= 3'b000;
      memory_array[5779] <= 3'b000;
      memory_array[5780] <= 3'b110;
      memory_array[5781] <= 3'b110;
      memory_array[5782] <= 3'b101;
      memory_array[5783] <= 3'b101;
      memory_array[5784] <= 3'b000;
      memory_array[5785] <= 3'b110;
      memory_array[5786] <= 3'b000;
      memory_array[5787] <= 3'b000;
      memory_array[5788] <= 3'b000;
      memory_array[5789] <= 3'b000;
      memory_array[5790] <= 3'b000;
      memory_array[5791] <= 3'b101;
      memory_array[5792] <= 3'b101;
      memory_array[5793] <= 3'b101;
      memory_array[5794] <= 3'b101;
      memory_array[5795] <= 3'b101;
      memory_array[5796] <= 3'b101;
      memory_array[5797] <= 3'b101;
      memory_array[5798] <= 3'b101;
      memory_array[5799] <= 3'b101;
      memory_array[5800] <= 3'b101;
      memory_array[5801] <= 3'b101;
      memory_array[5802] <= 3'b101;
      memory_array[5803] <= 3'b101;
      memory_array[5804] <= 3'b101;
      memory_array[5805] <= 3'b101;
      memory_array[5806] <= 3'b101;
      memory_array[5807] <= 3'b101;
      memory_array[5808] <= 3'b101;
      memory_array[5809] <= 3'b000;
      memory_array[5810] <= 3'b000;
      memory_array[5811] <= 3'b000;
      memory_array[5812] <= 3'b101;
      memory_array[5813] <= 3'b000;
      memory_array[5814] <= 3'b000;
      memory_array[5815] <= 3'b101;
      memory_array[5816] <= 3'b000;
      memory_array[5817] <= 3'b110;
      memory_array[5818] <= 3'b000;
      memory_array[5819] <= 3'b000;
      memory_array[5820] <= 3'b110;
      memory_array[5821] <= 3'b110;
      memory_array[5822] <= 3'b110;
      memory_array[5823] <= 3'b000;
      memory_array[5824] <= 3'b000;
      memory_array[5825] <= 3'b000;
      memory_array[5826] <= 3'b000;
      memory_array[5827] <= 3'b111;
      memory_array[5828] <= 3'b000;
      memory_array[5829] <= 3'b000;
      memory_array[5830] <= 3'b110;
      memory_array[5831] <= 3'b110;
      memory_array[5832] <= 3'b000;
      memory_array[5833] <= 3'b000;
      memory_array[5834] <= 3'b000;
      memory_array[5835] <= 3'b110;
      memory_array[5836] <= 3'b110;
      memory_array[5837] <= 3'b110;
      memory_array[5838] <= 3'b000;
      memory_array[5839] <= 3'b101;
      memory_array[5840] <= 3'b000;
      memory_array[5841] <= 3'b000;
      memory_array[5842] <= 3'b000;
      memory_array[5843] <= 3'b000;
      memory_array[5844] <= 3'b000;
      memory_array[5845] <= 3'b110;
      memory_array[5846] <= 3'b000;
      memory_array[5847] <= 3'b101;
      memory_array[5848] <= 3'b111;
      memory_array[5849] <= 3'b111;
      memory_array[5850] <= 3'b111;
      memory_array[5851] <= 3'b111;
      memory_array[5852] <= 3'b111;
      memory_array[5853] <= 3'b101;
      memory_array[5854] <= 3'b000;
      memory_array[5855] <= 3'b000;
      memory_array[5856] <= 3'b000;
      memory_array[5857] <= 3'b000;
      memory_array[5858] <= 3'b101;
      memory_array[5859] <= 3'b101;
      memory_array[5860] <= 3'b000;
      memory_array[5861] <= 3'b101;
      memory_array[5862] <= 3'b000;
      memory_array[5863] <= 3'b000;
      memory_array[5864] <= 3'b000;
      memory_array[5865] <= 3'b000;
      memory_array[5866] <= 3'b101;
      memory_array[5867] <= 3'b000;
      memory_array[5868] <= 3'b000;
      memory_array[5869] <= 3'b101;
      memory_array[5870] <= 3'b101;
      memory_array[5871] <= 3'b101;
      memory_array[5872] <= 3'b101;
      memory_array[5873] <= 3'b101;
      memory_array[5874] <= 3'b000;
      memory_array[5875] <= 3'b101;
      memory_array[5876] <= 3'b000;
      memory_array[5877] <= 3'b000;
      memory_array[5878] <= 3'b101;
      memory_array[5879] <= 3'b000;
      memory_array[5880] <= 3'b101;
      memory_array[5881] <= 3'b101;
      memory_array[5882] <= 3'b000;
      memory_array[5883] <= 3'b000;
      memory_array[5884] <= 3'b000;
      memory_array[5885] <= 3'b101;
      memory_array[5886] <= 3'b101;
      memory_array[5887] <= 3'b111;
      memory_array[5888] <= 3'b111;
      memory_array[5889] <= 3'b000;
      memory_array[5890] <= 3'b101;
      memory_array[5891] <= 3'b101;
      memory_array[5892] <= 3'b101;
      memory_array[5893] <= 3'b111;
      memory_array[5894] <= 3'b111;
      memory_array[5895] <= 3'b000;
      memory_array[5896] <= 3'b101;
      memory_array[5897] <= 3'b101;
      memory_array[5898] <= 3'b101;
      memory_array[5899] <= 3'b101;
      memory_array[5900] <= 3'b101;
      memory_array[5901] <= 3'b101;
      memory_array[5902] <= 3'b000;
      memory_array[5903] <= 3'b101;
      memory_array[5904] <= 3'b101;
      memory_array[5905] <= 3'b101;
      memory_array[5906] <= 3'b101;
      memory_array[5907] <= 3'b000;
      memory_array[5908] <= 3'b000;
      memory_array[5909] <= 3'b000;
      memory_array[5910] <= 3'b101;
      memory_array[5911] <= 3'b000;
      memory_array[5912] <= 3'b000;
      memory_array[5913] <= 3'b000;
      memory_array[5914] <= 3'b000;
      memory_array[5915] <= 3'b101;
      memory_array[5916] <= 3'b000;
      memory_array[5917] <= 3'b101;
      memory_array[5918] <= 3'b101;
      memory_array[5919] <= 3'b101;
      memory_array[5920] <= 3'b000;
      memory_array[5921] <= 3'b101;
      memory_array[5922] <= 3'b101;
      memory_array[5923] <= 3'b101;
      memory_array[5924] <= 3'b000;
      memory_array[5925] <= 3'b101;
      memory_array[5926] <= 3'b101;
      memory_array[5927] <= 3'b101;
      memory_array[5928] <= 3'b000;
      memory_array[5929] <= 3'b000;
      memory_array[5930] <= 3'b101;
      memory_array[5931] <= 3'b101;
      memory_array[5932] <= 3'b101;
      memory_array[5933] <= 3'b000;
      memory_array[5934] <= 3'b000;
      memory_array[5935] <= 3'b000;
      memory_array[5936] <= 3'b000;
      memory_array[5937] <= 3'b101;
      memory_array[5938] <= 3'b101;
      memory_array[5939] <= 3'b000;
      memory_array[5940] <= 3'b101;
      memory_array[5941] <= 3'b101;
      memory_array[5942] <= 3'b101;
      memory_array[5943] <= 3'b000;
      memory_array[5944] <= 3'b000;
      memory_array[5945] <= 3'b000;
      memory_array[5946] <= 3'b101;
      memory_array[5947] <= 3'b111;
      memory_array[5948] <= 3'b111;
      memory_array[5949] <= 3'b111;
      memory_array[5950] <= 3'b111;
      memory_array[5951] <= 3'b111;
      memory_array[5952] <= 3'b000;
      memory_array[5953] <= 3'b000;
      memory_array[5954] <= 3'b000;
      memory_array[5955] <= 3'b110;
      memory_array[5956] <= 3'b110;
      memory_array[5957] <= 3'b101;
      memory_array[5958] <= 3'b000;
      memory_array[5959] <= 3'b000;
      memory_array[5960] <= 3'b101;
      memory_array[5961] <= 3'b000;
      memory_array[5962] <= 3'b000;
      memory_array[5963] <= 3'b000;
      memory_array[5964] <= 3'b000;
      memory_array[5965] <= 3'b110;
      memory_array[5966] <= 3'b000;
      memory_array[5967] <= 3'b110;
      memory_array[5968] <= 3'b000;
      memory_array[5969] <= 3'b000;
      memory_array[5970] <= 3'b110;
      memory_array[5971] <= 3'b000;
      memory_array[5972] <= 3'b101;
      memory_array[5973] <= 3'b000;
      memory_array[5974] <= 3'b000;
      memory_array[5975] <= 3'b101;
      memory_array[5976] <= 3'b000;
      memory_array[5977] <= 3'b110;
      memory_array[5978] <= 3'b000;
      memory_array[5979] <= 3'b000;
      memory_array[5980] <= 3'b110;
      memory_array[5981] <= 3'b110;
      memory_array[5982] <= 3'b000;
      memory_array[5983] <= 3'b000;
      memory_array[5984] <= 3'b101;
      memory_array[5985] <= 3'b000;
      memory_array[5986] <= 3'b000;
      memory_array[5987] <= 3'b000;
      memory_array[5988] <= 3'b000;
      memory_array[5989] <= 3'b000;
      memory_array[5990] <= 3'b000;
      memory_array[5991] <= 3'b101;
      memory_array[5992] <= 3'b101;
      memory_array[5993] <= 3'b101;
      memory_array[5994] <= 3'b101;
      memory_array[5995] <= 3'b101;
      memory_array[5996] <= 3'b101;
      memory_array[5997] <= 3'b101;
      memory_array[5998] <= 3'b101;
      memory_array[5999] <= 3'b101;
      memory_array[6000] <= 3'b101;
      memory_array[6001] <= 3'b101;
      memory_array[6002] <= 3'b101;
      memory_array[6003] <= 3'b111;
      memory_array[6004] <= 3'b111;
      memory_array[6005] <= 3'b101;
      memory_array[6006] <= 3'b101;
      memory_array[6007] <= 3'b101;
      memory_array[6008] <= 3'b101;
      memory_array[6009] <= 3'b000;
      memory_array[6010] <= 3'b000;
      memory_array[6011] <= 3'b000;
      memory_array[6012] <= 3'b000;
      memory_array[6013] <= 3'b000;
      memory_array[6014] <= 3'b000;
      memory_array[6015] <= 3'b101;
      memory_array[6016] <= 3'b000;
      memory_array[6017] <= 3'b000;
      memory_array[6018] <= 3'b110;
      memory_array[6019] <= 3'b110;
      memory_array[6020] <= 3'b000;
      memory_array[6021] <= 3'b000;
      memory_array[6022] <= 3'b000;
      memory_array[6023] <= 3'b000;
      memory_array[6024] <= 3'b110;
      memory_array[6025] <= 3'b000;
      memory_array[6026] <= 3'b000;
      memory_array[6027] <= 3'b000;
      memory_array[6028] <= 3'b110;
      memory_array[6029] <= 3'b110;
      memory_array[6030] <= 3'b000;
      memory_array[6031] <= 3'b000;
      memory_array[6032] <= 3'b000;
      memory_array[6033] <= 3'b110;
      memory_array[6034] <= 3'b110;
      memory_array[6035] <= 3'b000;
      memory_array[6036] <= 3'b000;
      memory_array[6037] <= 3'b000;
      memory_array[6038] <= 3'b000;
      memory_array[6039] <= 3'b000;
      memory_array[6040] <= 3'b000;
      memory_array[6041] <= 3'b000;
      memory_array[6042] <= 3'b000;
      memory_array[6043] <= 3'b110;
      memory_array[6044] <= 3'b110;
      memory_array[6045] <= 3'b000;
      memory_array[6046] <= 3'b101;
      memory_array[6047] <= 3'b111;
      memory_array[6048] <= 3'b111;
      memory_array[6049] <= 3'b111;
      memory_array[6050] <= 3'b111;
      memory_array[6051] <= 3'b111;
      memory_array[6052] <= 3'b101;
      memory_array[6053] <= 3'b000;
      memory_array[6054] <= 3'b101;
      memory_array[6055] <= 3'b000;
      memory_array[6056] <= 3'b000;
      memory_array[6057] <= 3'b000;
      memory_array[6058] <= 3'b101;
      memory_array[6059] <= 3'b101;
      memory_array[6060] <= 3'b000;
      memory_array[6061] <= 3'b000;
      memory_array[6062] <= 3'b101;
      memory_array[6063] <= 3'b000;
      memory_array[6064] <= 3'b000;
      memory_array[6065] <= 3'b000;
      memory_array[6066] <= 3'b000;
      memory_array[6067] <= 3'b000;
      memory_array[6068] <= 3'b000;
      memory_array[6069] <= 3'b101;
      memory_array[6070] <= 3'b101;
      memory_array[6071] <= 3'b000;
      memory_array[6072] <= 3'b101;
      memory_array[6073] <= 3'b101;
      memory_array[6074] <= 3'b101;
      memory_array[6075] <= 3'b000;
      memory_array[6076] <= 3'b000;
      memory_array[6077] <= 3'b000;
      memory_array[6078] <= 3'b101;
      memory_array[6079] <= 3'b101;
      memory_array[6080] <= 3'b101;
      memory_array[6081] <= 3'b101;
      memory_array[6082] <= 3'b101;
      memory_array[6083] <= 3'b101;
      memory_array[6084] <= 3'b101;
      memory_array[6085] <= 3'b000;
      memory_array[6086] <= 3'b101;
      memory_array[6087] <= 3'b111;
      memory_array[6088] <= 3'b101;
      memory_array[6089] <= 3'b000;
      memory_array[6090] <= 3'b101;
      memory_array[6091] <= 3'b101;
      memory_array[6092] <= 3'b101;
      memory_array[6093] <= 3'b101;
      memory_array[6094] <= 3'b101;
      memory_array[6095] <= 3'b000;
      memory_array[6096] <= 3'b101;
      memory_array[6097] <= 3'b101;
      memory_array[6098] <= 3'b101;
      memory_array[6099] <= 3'b101;
      memory_array[6100] <= 3'b101;
      memory_array[6101] <= 3'b101;
      memory_array[6102] <= 3'b000;
      memory_array[6103] <= 3'b101;
      memory_array[6104] <= 3'b101;
      memory_array[6105] <= 3'b101;
      memory_array[6106] <= 3'b000;
      memory_array[6107] <= 3'b101;
      memory_array[6108] <= 3'b101;
      memory_array[6109] <= 3'b101;
      memory_array[6110] <= 3'b000;
      memory_array[6111] <= 3'b101;
      memory_array[6112] <= 3'b101;
      memory_array[6113] <= 3'b101;
      memory_array[6114] <= 3'b101;
      memory_array[6115] <= 3'b101;
      memory_array[6116] <= 3'b101;
      memory_array[6117] <= 3'b101;
      memory_array[6118] <= 3'b101;
      memory_array[6119] <= 3'b101;
      memory_array[6120] <= 3'b101;
      memory_array[6121] <= 3'b000;
      memory_array[6122] <= 3'b000;
      memory_array[6123] <= 3'b101;
      memory_array[6124] <= 3'b000;
      memory_array[6125] <= 3'b101;
      memory_array[6126] <= 3'b000;
      memory_array[6127] <= 3'b000;
      memory_array[6128] <= 3'b000;
      memory_array[6129] <= 3'b101;
      memory_array[6130] <= 3'b101;
      memory_array[6131] <= 3'b000;
      memory_array[6132] <= 3'b101;
      memory_array[6133] <= 3'b000;
      memory_array[6134] <= 3'b000;
      memory_array[6135] <= 3'b000;
      memory_array[6136] <= 3'b000;
      memory_array[6137] <= 3'b000;
      memory_array[6138] <= 3'b000;
      memory_array[6139] <= 3'b000;
      memory_array[6140] <= 3'b101;
      memory_array[6141] <= 3'b000;
      memory_array[6142] <= 3'b101;
      memory_array[6143] <= 3'b000;
      memory_array[6144] <= 3'b000;
      memory_array[6145] <= 3'b000;
      memory_array[6146] <= 3'b000;
      memory_array[6147] <= 3'b111;
      memory_array[6148] <= 3'b111;
      memory_array[6149] <= 3'b111;
      memory_array[6150] <= 3'b111;
      memory_array[6151] <= 3'b111;
      memory_array[6152] <= 3'b111;
      memory_array[6153] <= 3'b101;
      memory_array[6154] <= 3'b110;
      memory_array[6155] <= 3'b000;
      memory_array[6156] <= 3'b000;
      memory_array[6157] <= 3'b101;
      memory_array[6158] <= 3'b000;
      memory_array[6159] <= 3'b110;
      memory_array[6160] <= 3'b000;
      memory_array[6161] <= 3'b000;
      memory_array[6162] <= 3'b000;
      memory_array[6163] <= 3'b110;
      memory_array[6164] <= 3'b110;
      memory_array[6165] <= 3'b000;
      memory_array[6166] <= 3'b000;
      memory_array[6167] <= 3'b000;
      memory_array[6168] <= 3'b110;
      memory_array[6169] <= 3'b110;
      memory_array[6170] <= 3'b000;
      memory_array[6171] <= 3'b000;
      memory_array[6172] <= 3'b000;
      memory_array[6173] <= 3'b000;
      memory_array[6174] <= 3'b000;
      memory_array[6175] <= 3'b000;
      memory_array[6176] <= 3'b000;
      memory_array[6177] <= 3'b000;
      memory_array[6178] <= 3'b110;
      memory_array[6179] <= 3'b110;
      memory_array[6180] <= 3'b000;
      memory_array[6181] <= 3'b000;
      memory_array[6182] <= 3'b000;
      memory_array[6183] <= 3'b110;
      memory_array[6184] <= 3'b101;
      memory_array[6185] <= 3'b000;
      memory_array[6186] <= 3'b000;
      memory_array[6187] <= 3'b000;
      memory_array[6188] <= 3'b000;
      memory_array[6189] <= 3'b000;
      memory_array[6190] <= 3'b000;
      memory_array[6191] <= 3'b101;
      memory_array[6192] <= 3'b101;
      memory_array[6193] <= 3'b101;
      memory_array[6194] <= 3'b101;
      memory_array[6195] <= 3'b111;
      memory_array[6196] <= 3'b111;
      memory_array[6197] <= 3'b101;
      memory_array[6198] <= 3'b101;
      memory_array[6199] <= 3'b101;
      memory_array[6200] <= 3'b101;
      memory_array[6201] <= 3'b101;
      memory_array[6202] <= 3'b110;
      memory_array[6203] <= 3'b101;
      memory_array[6204] <= 3'b101;
      memory_array[6205] <= 3'b110;
      memory_array[6206] <= 3'b101;
      memory_array[6207] <= 3'b101;
      memory_array[6208] <= 3'b101;
      memory_array[6209] <= 3'b000;
      memory_array[6210] <= 3'b000;
      memory_array[6211] <= 3'b110;
      memory_array[6212] <= 3'b101;
      memory_array[6213] <= 3'b000;
      memory_array[6214] <= 3'b000;
      memory_array[6215] <= 3'b101;
      memory_array[6216] <= 3'b110;
      memory_array[6217] <= 3'b110;
      memory_array[6218] <= 3'b000;
      memory_array[6219] <= 3'b000;
      memory_array[6220] <= 3'b101;
      memory_array[6221] <= 3'b101;
      memory_array[6222] <= 3'b000;
      memory_array[6223] <= 3'b000;
      memory_array[6224] <= 3'b000;
      memory_array[6225] <= 3'b101;
      memory_array[6226] <= 3'b101;
      memory_array[6227] <= 3'b110;
      memory_array[6228] <= 3'b000;
      memory_array[6229] <= 3'b000;
      memory_array[6230] <= 3'b101;
      memory_array[6231] <= 3'b000;
      memory_array[6232] <= 3'b110;
      memory_array[6233] <= 3'b000;
      memory_array[6234] <= 3'b000;
      memory_array[6235] <= 3'b110;
      memory_array[6236] <= 3'b110;
      memory_array[6237] <= 3'b110;
      memory_array[6238] <= 3'b000;
      memory_array[6239] <= 3'b000;
      memory_array[6240] <= 3'b110;
      memory_array[6241] <= 3'b000;
      memory_array[6242] <= 3'b110;
      memory_array[6243] <= 3'b000;
      memory_array[6244] <= 3'b000;
      memory_array[6245] <= 3'b000;
      memory_array[6246] <= 3'b111;
      memory_array[6247] <= 3'b111;
      memory_array[6248] <= 3'b111;
      memory_array[6249] <= 3'b111;
      memory_array[6250] <= 3'b111;
      memory_array[6251] <= 3'b101;
      memory_array[6252] <= 3'b000;
      memory_array[6253] <= 3'b000;
      memory_array[6254] <= 3'b000;
      memory_array[6255] <= 3'b000;
      memory_array[6256] <= 3'b000;
      memory_array[6257] <= 3'b000;
      memory_array[6258] <= 3'b000;
      memory_array[6259] <= 3'b101;
      memory_array[6260] <= 3'b000;
      memory_array[6261] <= 3'b101;
      memory_array[6262] <= 3'b101;
      memory_array[6263] <= 3'b000;
      memory_array[6264] <= 3'b101;
      memory_array[6265] <= 3'b000;
      memory_array[6266] <= 3'b000;
      memory_array[6267] <= 3'b000;
      memory_array[6268] <= 3'b000;
      memory_array[6269] <= 3'b000;
      memory_array[6270] <= 3'b101;
      memory_array[6271] <= 3'b101;
      memory_array[6272] <= 3'b000;
      memory_array[6273] <= 3'b000;
      memory_array[6274] <= 3'b000;
      memory_array[6275] <= 3'b101;
      memory_array[6276] <= 3'b000;
      memory_array[6277] <= 3'b101;
      memory_array[6278] <= 3'b101;
      memory_array[6279] <= 3'b101;
      memory_array[6280] <= 3'b101;
      memory_array[6281] <= 3'b000;
      memory_array[6282] <= 3'b000;
      memory_array[6283] <= 3'b000;
      memory_array[6284] <= 3'b101;
      memory_array[6285] <= 3'b000;
      memory_array[6286] <= 3'b101;
      memory_array[6287] <= 3'b101;
      memory_array[6288] <= 3'b000;
      memory_array[6289] <= 3'b000;
      memory_array[6290] <= 3'b101;
      memory_array[6291] <= 3'b000;
      memory_array[6292] <= 3'b101;
      memory_array[6293] <= 3'b000;
      memory_array[6294] <= 3'b000;
      memory_array[6295] <= 3'b000;
      memory_array[6296] <= 3'b000;
      memory_array[6297] <= 3'b000;
      memory_array[6298] <= 3'b101;
      memory_array[6299] <= 3'b101;
      memory_array[6300] <= 3'b101;
      memory_array[6301] <= 3'b101;
      memory_array[6302] <= 3'b101;
      memory_array[6303] <= 3'b101;
      memory_array[6304] <= 3'b000;
      memory_array[6305] <= 3'b101;
      memory_array[6306] <= 3'b101;
      memory_array[6307] <= 3'b101;
      memory_array[6308] <= 3'b101;
      memory_array[6309] <= 3'b101;
      memory_array[6310] <= 3'b101;
      memory_array[6311] <= 3'b101;
      memory_array[6312] <= 3'b000;
      memory_array[6313] <= 3'b101;
      memory_array[6314] <= 3'b000;
      memory_array[6315] <= 3'b101;
      memory_array[6316] <= 3'b000;
      memory_array[6317] <= 3'b101;
      memory_array[6318] <= 3'b000;
      memory_array[6319] <= 3'b101;
      memory_array[6320] <= 3'b101;
      memory_array[6321] <= 3'b101;
      memory_array[6322] <= 3'b101;
      memory_array[6323] <= 3'b000;
      memory_array[6324] <= 3'b000;
      memory_array[6325] <= 3'b000;
      memory_array[6326] <= 3'b000;
      memory_array[6327] <= 3'b101;
      memory_array[6328] <= 3'b101;
      memory_array[6329] <= 3'b101;
      memory_array[6330] <= 3'b101;
      memory_array[6331] <= 3'b000;
      memory_array[6332] <= 3'b101;
      memory_array[6333] <= 3'b000;
      memory_array[6334] <= 3'b000;
      memory_array[6335] <= 3'b101;
      memory_array[6336] <= 3'b000;
      memory_array[6337] <= 3'b000;
      memory_array[6338] <= 3'b000;
      memory_array[6339] <= 3'b000;
      memory_array[6340] <= 3'b101;
      memory_array[6341] <= 3'b000;
      memory_array[6342] <= 3'b101;
      memory_array[6343] <= 3'b000;
      memory_array[6344] <= 3'b000;
      memory_array[6345] <= 3'b000;
      memory_array[6346] <= 3'b101;
      memory_array[6347] <= 3'b101;
      memory_array[6348] <= 3'b101;
      memory_array[6349] <= 3'b111;
      memory_array[6350] <= 3'b111;
      memory_array[6351] <= 3'b111;
      memory_array[6352] <= 3'b111;
      memory_array[6353] <= 3'b111;
      memory_array[6354] <= 3'b000;
      memory_array[6355] <= 3'b110;
      memory_array[6356] <= 3'b110;
      memory_array[6357] <= 3'b110;
      memory_array[6358] <= 3'b000;
      memory_array[6359] <= 3'b000;
      memory_array[6360] <= 3'b000;
      memory_array[6361] <= 3'b000;
      memory_array[6362] <= 3'b110;
      memory_array[6363] <= 3'b000;
      memory_array[6364] <= 3'b000;
      memory_array[6365] <= 3'b110;
      memory_array[6366] <= 3'b110;
      memory_array[6367] <= 3'b000;
      memory_array[6368] <= 3'b000;
      memory_array[6369] <= 3'b101;
      memory_array[6370] <= 3'b000;
      memory_array[6371] <= 3'b110;
      memory_array[6372] <= 3'b000;
      memory_array[6373] <= 3'b101;
      memory_array[6374] <= 3'b101;
      memory_array[6375] <= 3'b000;
      memory_array[6376] <= 3'b110;
      memory_array[6377] <= 3'b101;
      memory_array[6378] <= 3'b101;
      memory_array[6379] <= 3'b000;
      memory_array[6380] <= 3'b000;
      memory_array[6381] <= 3'b110;
      memory_array[6382] <= 3'b110;
      memory_array[6383] <= 3'b000;
      memory_array[6384] <= 3'b101;
      memory_array[6385] <= 3'b000;
      memory_array[6386] <= 3'b000;
      memory_array[6387] <= 3'b000;
      memory_array[6388] <= 3'b000;
      memory_array[6389] <= 3'b000;
      memory_array[6390] <= 3'b000;
      memory_array[6391] <= 3'b101;
      memory_array[6392] <= 3'b101;
      memory_array[6393] <= 3'b101;
      memory_array[6394] <= 3'b000;
      memory_array[6395] <= 3'b101;
      memory_array[6396] <= 3'b101;
      memory_array[6397] <= 3'b110;
      memory_array[6398] <= 3'b101;
      memory_array[6399] <= 3'b101;
      memory_array[6400] <= 3'b101;
      memory_array[6401] <= 3'b110;
      memory_array[6402] <= 3'b110;
      memory_array[6403] <= 3'b000;
      memory_array[6404] <= 3'b000;
      memory_array[6405] <= 3'b110;
      memory_array[6406] <= 3'b110;
      memory_array[6407] <= 3'b101;
      memory_array[6408] <= 3'b101;
      memory_array[6409] <= 3'b000;
      memory_array[6410] <= 3'b000;
      memory_array[6411] <= 3'b110;
      memory_array[6412] <= 3'b000;
      memory_array[6413] <= 3'b000;
      memory_array[6414] <= 3'b000;
      memory_array[6415] <= 3'b000;
      memory_array[6416] <= 3'b000;
      memory_array[6417] <= 3'b110;
      memory_array[6418] <= 3'b000;
      memory_array[6419] <= 3'b000;
      memory_array[6420] <= 3'b101;
      memory_array[6421] <= 3'b000;
      memory_array[6422] <= 3'b101;
      memory_array[6423] <= 3'b000;
      memory_array[6424] <= 3'b101;
      memory_array[6425] <= 3'b000;
      memory_array[6426] <= 3'b000;
      memory_array[6427] <= 3'b000;
      memory_array[6428] <= 3'b000;
      memory_array[6429] <= 3'b000;
      memory_array[6430] <= 3'b000;
      memory_array[6431] <= 3'b000;
      memory_array[6432] <= 3'b000;
      memory_array[6433] <= 3'b000;
      memory_array[6434] <= 3'b000;
      memory_array[6435] <= 3'b110;
      memory_array[6436] <= 3'b110;
      memory_array[6437] <= 3'b000;
      memory_array[6438] <= 3'b101;
      memory_array[6439] <= 3'b000;
      memory_array[6440] <= 3'b110;
      memory_array[6441] <= 3'b110;
      memory_array[6442] <= 3'b110;
      memory_array[6443] <= 3'b000;
      memory_array[6444] <= 3'b111;
      memory_array[6445] <= 3'b111;
      memory_array[6446] <= 3'b111;
      memory_array[6447] <= 3'b111;
      memory_array[6448] <= 3'b111;
      memory_array[6449] <= 3'b101;
      memory_array[6450] <= 3'b101;
      memory_array[6451] <= 3'b101;
      memory_array[6452] <= 3'b000;
      memory_array[6453] <= 3'b101;
      memory_array[6454] <= 3'b000;
      memory_array[6455] <= 3'b000;
      memory_array[6456] <= 3'b101;
      memory_array[6457] <= 3'b101;
      memory_array[6458] <= 3'b000;
      memory_array[6459] <= 3'b101;
      memory_array[6460] <= 3'b101;
      memory_array[6461] <= 3'b000;
      memory_array[6462] <= 3'b101;
      memory_array[6463] <= 3'b101;
      memory_array[6464] <= 3'b101;
      memory_array[6465] <= 3'b101;
      memory_array[6466] <= 3'b101;
      memory_array[6467] <= 3'b000;
      memory_array[6468] <= 3'b000;
      memory_array[6469] <= 3'b101;
      memory_array[6470] <= 3'b101;
      memory_array[6471] <= 3'b000;
      memory_array[6472] <= 3'b000;
      memory_array[6473] <= 3'b000;
      memory_array[6474] <= 3'b101;
      memory_array[6475] <= 3'b101;
      memory_array[6476] <= 3'b101;
      memory_array[6477] <= 3'b000;
      memory_array[6478] <= 3'b101;
      memory_array[6479] <= 3'b101;
      memory_array[6480] <= 3'b101;
      memory_array[6481] <= 3'b000;
      memory_array[6482] <= 3'b101;
      memory_array[6483] <= 3'b000;
      memory_array[6484] <= 3'b101;
      memory_array[6485] <= 3'b000;
      memory_array[6486] <= 3'b101;
      memory_array[6487] <= 3'b101;
      memory_array[6488] <= 3'b000;
      memory_array[6489] <= 3'b101;
      memory_array[6490] <= 3'b000;
      memory_array[6491] <= 3'b000;
      memory_array[6492] <= 3'b101;
      memory_array[6493] <= 3'b101;
      memory_array[6494] <= 3'b000;
      memory_array[6495] <= 3'b000;
      memory_array[6496] <= 3'b101;
      memory_array[6497] <= 3'b101;
      memory_array[6498] <= 3'b000;
      memory_array[6499] <= 3'b000;
      memory_array[6500] <= 3'b000;
      memory_array[6501] <= 3'b101;
      memory_array[6502] <= 3'b101;
      memory_array[6503] <= 3'b101;
      memory_array[6504] <= 3'b101;
      memory_array[6505] <= 3'b000;
      memory_array[6506] <= 3'b101;
      memory_array[6507] <= 3'b000;
      memory_array[6508] <= 3'b000;
      memory_array[6509] <= 3'b101;
      memory_array[6510] <= 3'b101;
      memory_array[6511] <= 3'b000;
      memory_array[6512] <= 3'b101;
      memory_array[6513] <= 3'b101;
      memory_array[6514] <= 3'b000;
      memory_array[6515] <= 3'b101;
      memory_array[6516] <= 3'b000;
      memory_array[6517] <= 3'b101;
      memory_array[6518] <= 3'b000;
      memory_array[6519] <= 3'b101;
      memory_array[6520] <= 3'b101;
      memory_array[6521] <= 3'b101;
      memory_array[6522] <= 3'b101;
      memory_array[6523] <= 3'b101;
      memory_array[6524] <= 3'b101;
      memory_array[6525] <= 3'b101;
      memory_array[6526] <= 3'b000;
      memory_array[6527] <= 3'b101;
      memory_array[6528] <= 3'b000;
      memory_array[6529] <= 3'b101;
      memory_array[6530] <= 3'b101;
      memory_array[6531] <= 3'b000;
      memory_array[6532] <= 3'b000;
      memory_array[6533] <= 3'b101;
      memory_array[6534] <= 3'b101;
      memory_array[6535] <= 3'b101;
      memory_array[6536] <= 3'b101;
      memory_array[6537] <= 3'b000;
      memory_array[6538] <= 3'b000;
      memory_array[6539] <= 3'b101;
      memory_array[6540] <= 3'b101;
      memory_array[6541] <= 3'b000;
      memory_array[6542] <= 3'b000;
      memory_array[6543] <= 3'b101;
      memory_array[6544] <= 3'b000;
      memory_array[6545] <= 3'b000;
      memory_array[6546] <= 3'b101;
      memory_array[6547] <= 3'b101;
      memory_array[6548] <= 3'b000;
      memory_array[6549] <= 3'b101;
      memory_array[6550] <= 3'b101;
      memory_array[6551] <= 3'b111;
      memory_array[6552] <= 3'b111;
      memory_array[6553] <= 3'b111;
      memory_array[6554] <= 3'b111;
      memory_array[6555] <= 3'b111;
      memory_array[6556] <= 3'b000;
      memory_array[6557] <= 3'b110;
      memory_array[6558] <= 3'b000;
      memory_array[6559] <= 3'b000;
      memory_array[6560] <= 3'b110;
      memory_array[6561] <= 3'b101;
      memory_array[6562] <= 3'b110;
      memory_array[6563] <= 3'b000;
      memory_array[6564] <= 3'b000;
      memory_array[6565] <= 3'b110;
      memory_array[6566] <= 3'b110;
      memory_array[6567] <= 3'b101;
      memory_array[6568] <= 3'b000;
      memory_array[6569] <= 3'b000;
      memory_array[6570] <= 3'b000;
      memory_array[6571] <= 3'b000;
      memory_array[6572] <= 3'b101;
      memory_array[6573] <= 3'b000;
      memory_array[6574] <= 3'b000;
      memory_array[6575] <= 3'b101;
      memory_array[6576] <= 3'b000;
      memory_array[6577] <= 3'b000;
      memory_array[6578] <= 3'b000;
      memory_array[6579] <= 3'b101;
      memory_array[6580] <= 3'b101;
      memory_array[6581] <= 3'b110;
      memory_array[6582] <= 3'b110;
      memory_array[6583] <= 3'b000;
      memory_array[6584] <= 3'b000;
      memory_array[6585] <= 3'b110;
      memory_array[6586] <= 3'b000;
      memory_array[6587] <= 3'b000;
      memory_array[6588] <= 3'b000;
      memory_array[6589] <= 3'b000;
      memory_array[6590] <= 3'b000;
      memory_array[6591] <= 3'b101;
      memory_array[6592] <= 3'b110;
      memory_array[6593] <= 3'b000;
      memory_array[6594] <= 3'b000;
      memory_array[6595] <= 3'b110;
      memory_array[6596] <= 3'b110;
      memory_array[6597] <= 3'b110;
      memory_array[6598] <= 3'b000;
      memory_array[6599] <= 3'b101;
      memory_array[6600] <= 3'b000;
      memory_array[6601] <= 3'b000;
      memory_array[6602] <= 3'b000;
      memory_array[6603] <= 3'b110;
      memory_array[6604] <= 3'b110;
      memory_array[6605] <= 3'b000;
      memory_array[6606] <= 3'b000;
      memory_array[6607] <= 3'b000;
      memory_array[6608] <= 3'b101;
      memory_array[6609] <= 3'b000;
      memory_array[6610] <= 3'b000;
      memory_array[6611] <= 3'b000;
      memory_array[6612] <= 3'b000;
      memory_array[6613] <= 3'b000;
      memory_array[6614] <= 3'b110;
      memory_array[6615] <= 3'b000;
      memory_array[6616] <= 3'b000;
      memory_array[6617] <= 3'b000;
      memory_array[6618] <= 3'b110;
      memory_array[6619] <= 3'b101;
      memory_array[6620] <= 3'b000;
      memory_array[6621] <= 3'b000;
      memory_array[6622] <= 3'b101;
      memory_array[6623] <= 3'b101;
      memory_array[6624] <= 3'b101;
      memory_array[6625] <= 3'b000;
      memory_array[6626] <= 3'b000;
      memory_array[6627] <= 3'b000;
      memory_array[6628] <= 3'b000;
      memory_array[6629] <= 3'b000;
      memory_array[6630] <= 3'b000;
      memory_array[6631] <= 3'b000;
      memory_array[6632] <= 3'b000;
      memory_array[6633] <= 3'b110;
      memory_array[6634] <= 3'b110;
      memory_array[6635] <= 3'b000;
      memory_array[6636] <= 3'b000;
      memory_array[6637] <= 3'b000;
      memory_array[6638] <= 3'b110;
      memory_array[6639] <= 3'b110;
      memory_array[6640] <= 3'b000;
      memory_array[6641] <= 3'b000;
      memory_array[6642] <= 3'b000;
      memory_array[6643] <= 3'b101;
      memory_array[6644] <= 3'b111;
      memory_array[6645] <= 3'b111;
      memory_array[6646] <= 3'b111;
      memory_array[6647] <= 3'b111;
      memory_array[6648] <= 3'b111;
      memory_array[6649] <= 3'b000;
      memory_array[6650] <= 3'b000;
      memory_array[6651] <= 3'b000;
      memory_array[6652] <= 3'b000;
      memory_array[6653] <= 3'b000;
      memory_array[6654] <= 3'b101;
      memory_array[6655] <= 3'b000;
      memory_array[6656] <= 3'b101;
      memory_array[6657] <= 3'b000;
      memory_array[6658] <= 3'b000;
      memory_array[6659] <= 3'b101;
      memory_array[6660] <= 3'b000;
      memory_array[6661] <= 3'b101;
      memory_array[6662] <= 3'b101;
      memory_array[6663] <= 3'b101;
      memory_array[6664] <= 3'b000;
      memory_array[6665] <= 3'b101;
      memory_array[6666] <= 3'b101;
      memory_array[6667] <= 3'b000;
      memory_array[6668] <= 3'b101;
      memory_array[6669] <= 3'b101;
      memory_array[6670] <= 3'b101;
      memory_array[6671] <= 3'b000;
      memory_array[6672] <= 3'b101;
      memory_array[6673] <= 3'b101;
      memory_array[6674] <= 3'b101;
      memory_array[6675] <= 3'b101;
      memory_array[6676] <= 3'b000;
      memory_array[6677] <= 3'b000;
      memory_array[6678] <= 3'b101;
      memory_array[6679] <= 3'b101;
      memory_array[6680] <= 3'b000;
      memory_array[6681] <= 3'b000;
      memory_array[6682] <= 3'b101;
      memory_array[6683] <= 3'b101;
      memory_array[6684] <= 3'b101;
      memory_array[6685] <= 3'b000;
      memory_array[6686] <= 3'b101;
      memory_array[6687] <= 3'b111;
      memory_array[6688] <= 3'b000;
      memory_array[6689] <= 3'b101;
      memory_array[6690] <= 3'b000;
      memory_array[6691] <= 3'b000;
      memory_array[6692] <= 3'b101;
      memory_array[6693] <= 3'b111;
      memory_array[6694] <= 3'b000;
      memory_array[6695] <= 3'b000;
      memory_array[6696] <= 3'b000;
      memory_array[6697] <= 3'b101;
      memory_array[6698] <= 3'b000;
      memory_array[6699] <= 3'b101;
      memory_array[6700] <= 3'b101;
      memory_array[6701] <= 3'b101;
      memory_array[6702] <= 3'b000;
      memory_array[6703] <= 3'b000;
      memory_array[6704] <= 3'b101;
      memory_array[6705] <= 3'b101;
      memory_array[6706] <= 3'b101;
      memory_array[6707] <= 3'b101;
      memory_array[6708] <= 3'b000;
      memory_array[6709] <= 3'b000;
      memory_array[6710] <= 3'b101;
      memory_array[6711] <= 3'b000;
      memory_array[6712] <= 3'b101;
      memory_array[6713] <= 3'b101;
      memory_array[6714] <= 3'b000;
      memory_array[6715] <= 3'b101;
      memory_array[6716] <= 3'b000;
      memory_array[6717] <= 3'b101;
      memory_array[6718] <= 3'b101;
      memory_array[6719] <= 3'b000;
      memory_array[6720] <= 3'b101;
      memory_array[6721] <= 3'b000;
      memory_array[6722] <= 3'b000;
      memory_array[6723] <= 3'b000;
      memory_array[6724] <= 3'b101;
      memory_array[6725] <= 3'b000;
      memory_array[6726] <= 3'b101;
      memory_array[6727] <= 3'b101;
      memory_array[6728] <= 3'b101;
      memory_array[6729] <= 3'b101;
      memory_array[6730] <= 3'b101;
      memory_array[6731] <= 3'b101;
      memory_array[6732] <= 3'b000;
      memory_array[6733] <= 3'b101;
      memory_array[6734] <= 3'b101;
      memory_array[6735] <= 3'b000;
      memory_array[6736] <= 3'b101;
      memory_array[6737] <= 3'b000;
      memory_array[6738] <= 3'b101;
      memory_array[6739] <= 3'b000;
      memory_array[6740] <= 3'b101;
      memory_array[6741] <= 3'b000;
      memory_array[6742] <= 3'b000;
      memory_array[6743] <= 3'b101;
      memory_array[6744] <= 3'b000;
      memory_array[6745] <= 3'b101;
      memory_array[6746] <= 3'b000;
      memory_array[6747] <= 3'b101;
      memory_array[6748] <= 3'b000;
      memory_array[6749] <= 3'b000;
      memory_array[6750] <= 3'b000;
      memory_array[6751] <= 3'b111;
      memory_array[6752] <= 3'b111;
      memory_array[6753] <= 3'b111;
      memory_array[6754] <= 3'b111;
      memory_array[6755] <= 3'b111;
      memory_array[6756] <= 3'b101;
      memory_array[6757] <= 3'b000;
      memory_array[6758] <= 3'b110;
      memory_array[6759] <= 3'b110;
      memory_array[6760] <= 3'b000;
      memory_array[6761] <= 3'b000;
      memory_array[6762] <= 3'b000;
      memory_array[6763] <= 3'b110;
      memory_array[6764] <= 3'b110;
      memory_array[6765] <= 3'b000;
      memory_array[6766] <= 3'b000;
      memory_array[6767] <= 3'b000;
      memory_array[6768] <= 3'b000;
      memory_array[6769] <= 3'b110;
      memory_array[6770] <= 3'b000;
      memory_array[6771] <= 3'b000;
      memory_array[6772] <= 3'b000;
      memory_array[6773] <= 3'b000;
      memory_array[6774] <= 3'b000;
      memory_array[6775] <= 3'b000;
      memory_array[6776] <= 3'b000;
      memory_array[6777] <= 3'b000;
      memory_array[6778] <= 3'b110;
      memory_array[6779] <= 3'b101;
      memory_array[6780] <= 3'b101;
      memory_array[6781] <= 3'b000;
      memory_array[6782] <= 3'b000;
      memory_array[6783] <= 3'b110;
      memory_array[6784] <= 3'b000;
      memory_array[6785] <= 3'b000;
      memory_array[6786] <= 3'b000;
      memory_array[6787] <= 3'b000;
      memory_array[6788] <= 3'b110;
      memory_array[6789] <= 3'b000;
      memory_array[6790] <= 3'b000;
      memory_array[6791] <= 3'b101;
      memory_array[6792] <= 3'b000;
      memory_array[6793] <= 3'b110;
      memory_array[6794] <= 3'b110;
      memory_array[6795] <= 3'b000;
      memory_array[6796] <= 3'b000;
      memory_array[6797] <= 3'b000;
      memory_array[6798] <= 3'b110;
      memory_array[6799] <= 3'b110;
      memory_array[6800] <= 3'b101;
      memory_array[6801] <= 3'b101;
      memory_array[6802] <= 3'b101;
      memory_array[6803] <= 3'b101;
      memory_array[6804] <= 3'b101;
      memory_array[6805] <= 3'b101;
      memory_array[6806] <= 3'b101;
      memory_array[6807] <= 3'b101;
      memory_array[6808] <= 3'b101;
      memory_array[6809] <= 3'b000;
      memory_array[6810] <= 3'b000;
      memory_array[6811] <= 3'b000;
      memory_array[6812] <= 3'b101;
      memory_array[6813] <= 3'b000;
      memory_array[6814] <= 3'b101;
      memory_array[6815] <= 3'b101;
      memory_array[6816] <= 3'b000;
      memory_array[6817] <= 3'b000;
      memory_array[6818] <= 3'b110;
      memory_array[6819] <= 3'b110;
      memory_array[6820] <= 3'b000;
      memory_array[6821] <= 3'b000;
      memory_array[6822] <= 3'b101;
      memory_array[6823] <= 3'b101;
      memory_array[6824] <= 3'b110;
      memory_array[6825] <= 3'b000;
      memory_array[6826] <= 3'b000;
      memory_array[6827] <= 3'b000;
      memory_array[6828] <= 3'b000;
      memory_array[6829] <= 3'b101;
      memory_array[6830] <= 3'b000;
      memory_array[6831] <= 3'b000;
      memory_array[6832] <= 3'b101;
      memory_array[6833] <= 3'b101;
      memory_array[6834] <= 3'b000;
      memory_array[6835] <= 3'b000;
      memory_array[6836] <= 3'b000;
      memory_array[6837] <= 3'b000;
      memory_array[6838] <= 3'b110;
      memory_array[6839] <= 3'b111;
      memory_array[6840] <= 3'b000;
      memory_array[6841] <= 3'b000;
      memory_array[6842] <= 3'b111;
      memory_array[6843] <= 3'b111;
      memory_array[6844] <= 3'b111;
      memory_array[6845] <= 3'b111;
      memory_array[6846] <= 3'b111;
      memory_array[6847] <= 3'b101;
      memory_array[6848] <= 3'b000;
      memory_array[6849] <= 3'b101;
      memory_array[6850] <= 3'b101;
      memory_array[6851] <= 3'b000;
      memory_array[6852] <= 3'b000;
      memory_array[6853] <= 3'b000;
      memory_array[6854] <= 3'b101;
      memory_array[6855] <= 3'b000;
      memory_array[6856] <= 3'b000;
      memory_array[6857] <= 3'b000;
      memory_array[6858] <= 3'b101;
      memory_array[6859] <= 3'b000;
      memory_array[6860] <= 3'b101;
      memory_array[6861] <= 3'b101;
      memory_array[6862] <= 3'b101;
      memory_array[6863] <= 3'b000;
      memory_array[6864] <= 3'b101;
      memory_array[6865] <= 3'b101;
      memory_array[6866] <= 3'b101;
      memory_array[6867] <= 3'b101;
      memory_array[6868] <= 3'b101;
      memory_array[6869] <= 3'b101;
      memory_array[6870] <= 3'b101;
      memory_array[6871] <= 3'b101;
      memory_array[6872] <= 3'b101;
      memory_array[6873] <= 3'b000;
      memory_array[6874] <= 3'b101;
      memory_array[6875] <= 3'b000;
      memory_array[6876] <= 3'b101;
      memory_array[6877] <= 3'b101;
      memory_array[6878] <= 3'b000;
      memory_array[6879] <= 3'b101;
      memory_array[6880] <= 3'b101;
      memory_array[6881] <= 3'b101;
      memory_array[6882] <= 3'b000;
      memory_array[6883] <= 3'b000;
      memory_array[6884] <= 3'b101;
      memory_array[6885] <= 3'b000;
      memory_array[6886] <= 3'b111;
      memory_array[6887] <= 3'b111;
      memory_array[6888] <= 3'b111;
      memory_array[6889] <= 3'b000;
      memory_array[6890] <= 3'b000;
      memory_array[6891] <= 3'b101;
      memory_array[6892] <= 3'b111;
      memory_array[6893] <= 3'b111;
      memory_array[6894] <= 3'b111;
      memory_array[6895] <= 3'b111;
      memory_array[6896] <= 3'b101;
      memory_array[6897] <= 3'b101;
      memory_array[6898] <= 3'b000;
      memory_array[6899] <= 3'b101;
      memory_array[6900] <= 3'b000;
      memory_array[6901] <= 3'b101;
      memory_array[6902] <= 3'b000;
      memory_array[6903] <= 3'b000;
      memory_array[6904] <= 3'b101;
      memory_array[6905] <= 3'b000;
      memory_array[6906] <= 3'b101;
      memory_array[6907] <= 3'b101;
      memory_array[6908] <= 3'b000;
      memory_array[6909] <= 3'b101;
      memory_array[6910] <= 3'b101;
      memory_array[6911] <= 3'b000;
      memory_array[6912] <= 3'b000;
      memory_array[6913] <= 3'b000;
      memory_array[6914] <= 3'b000;
      memory_array[6915] <= 3'b101;
      memory_array[6916] <= 3'b000;
      memory_array[6917] <= 3'b101;
      memory_array[6918] <= 3'b101;
      memory_array[6919] <= 3'b101;
      memory_array[6920] <= 3'b101;
      memory_array[6921] <= 3'b000;
      memory_array[6922] <= 3'b101;
      memory_array[6923] <= 3'b101;
      memory_array[6924] <= 3'b000;
      memory_array[6925] <= 3'b101;
      memory_array[6926] <= 3'b000;
      memory_array[6927] <= 3'b101;
      memory_array[6928] <= 3'b101;
      memory_array[6929] <= 3'b101;
      memory_array[6930] <= 3'b101;
      memory_array[6931] <= 3'b101;
      memory_array[6932] <= 3'b101;
      memory_array[6933] <= 3'b101;
      memory_array[6934] <= 3'b101;
      memory_array[6935] <= 3'b101;
      memory_array[6936] <= 3'b000;
      memory_array[6937] <= 3'b000;
      memory_array[6938] <= 3'b101;
      memory_array[6939] <= 3'b101;
      memory_array[6940] <= 3'b000;
      memory_array[6941] <= 3'b101;
      memory_array[6942] <= 3'b101;
      memory_array[6943] <= 3'b000;
      memory_array[6944] <= 3'b000;
      memory_array[6945] <= 3'b101;
      memory_array[6946] <= 3'b000;
      memory_array[6947] <= 3'b000;
      memory_array[6948] <= 3'b000;
      memory_array[6949] <= 3'b101;
      memory_array[6950] <= 3'b000;
      memory_array[6951] <= 3'b000;
      memory_array[6952] <= 3'b101;
      memory_array[6953] <= 3'b111;
      memory_array[6954] <= 3'b111;
      memory_array[6955] <= 3'b111;
      memory_array[6956] <= 3'b111;
      memory_array[6957] <= 3'b101;
      memory_array[6958] <= 3'b000;
      memory_array[6959] <= 3'b000;
      memory_array[6960] <= 3'b111;
      memory_array[6961] <= 3'b000;
      memory_array[6962] <= 3'b101;
      memory_array[6963] <= 3'b000;
      memory_array[6964] <= 3'b110;
      memory_array[6965] <= 3'b000;
      memory_array[6966] <= 3'b101;
      memory_array[6967] <= 3'b000;
      memory_array[6968] <= 3'b110;
      memory_array[6969] <= 3'b000;
      memory_array[6970] <= 3'b101;
      memory_array[6971] <= 3'b000;
      memory_array[6972] <= 3'b000;
      memory_array[6973] <= 3'b110;
      memory_array[6974] <= 3'b110;
      memory_array[6975] <= 3'b000;
      memory_array[6976] <= 3'b000;
      memory_array[6977] <= 3'b101;
      memory_array[6978] <= 3'b000;
      memory_array[6979] <= 3'b110;
      memory_array[6980] <= 3'b000;
      memory_array[6981] <= 3'b000;
      memory_array[6982] <= 3'b000;
      memory_array[6983] <= 3'b110;
      memory_array[6984] <= 3'b101;
      memory_array[6985] <= 3'b101;
      memory_array[6986] <= 3'b000;
      memory_array[6987] <= 3'b101;
      memory_array[6988] <= 3'b000;
      memory_array[6989] <= 3'b000;
      memory_array[6990] <= 3'b000;
      memory_array[6991] <= 3'b101;
      memory_array[6992] <= 3'b101;
      memory_array[6993] <= 3'b101;
      memory_array[6994] <= 3'b101;
      memory_array[6995] <= 3'b101;
      memory_array[6996] <= 3'b101;
      memory_array[6997] <= 3'b101;
      memory_array[6998] <= 3'b101;
      memory_array[6999] <= 3'b101;
      memory_array[7000] <= 3'b101;
      memory_array[7001] <= 3'b101;
      memory_array[7002] <= 3'b101;
      memory_array[7003] <= 3'b101;
      memory_array[7004] <= 3'b101;
      memory_array[7005] <= 3'b101;
      memory_array[7006] <= 3'b101;
      memory_array[7007] <= 3'b101;
      memory_array[7008] <= 3'b101;
      memory_array[7009] <= 3'b000;
      memory_array[7010] <= 3'b000;
      memory_array[7011] <= 3'b000;
      memory_array[7012] <= 3'b101;
      memory_array[7013] <= 3'b000;
      memory_array[7014] <= 3'b101;
      memory_array[7015] <= 3'b101;
      memory_array[7016] <= 3'b000;
      memory_array[7017] <= 3'b000;
      memory_array[7018] <= 3'b110;
      memory_array[7019] <= 3'b110;
      memory_array[7020] <= 3'b000;
      memory_array[7021] <= 3'b000;
      memory_array[7022] <= 3'b101;
      memory_array[7023] <= 3'b101;
      memory_array[7024] <= 3'b110;
      memory_array[7025] <= 3'b000;
      memory_array[7026] <= 3'b000;
      memory_array[7027] <= 3'b000;
      memory_array[7028] <= 3'b000;
      memory_array[7029] <= 3'b101;
      memory_array[7030] <= 3'b000;
      memory_array[7031] <= 3'b000;
      memory_array[7032] <= 3'b101;
      memory_array[7033] <= 3'b101;
      memory_array[7034] <= 3'b000;
      memory_array[7035] <= 3'b000;
      memory_array[7036] <= 3'b000;
      memory_array[7037] <= 3'b000;
      memory_array[7038] <= 3'b110;
      memory_array[7039] <= 3'b111;
      memory_array[7040] <= 3'b000;
      memory_array[7041] <= 3'b000;
      memory_array[7042] <= 3'b111;
      memory_array[7043] <= 3'b111;
      memory_array[7044] <= 3'b111;
      memory_array[7045] <= 3'b111;
      memory_array[7046] <= 3'b111;
      memory_array[7047] <= 3'b101;
      memory_array[7048] <= 3'b000;
      memory_array[7049] <= 3'b101;
      memory_array[7050] <= 3'b101;
      memory_array[7051] <= 3'b000;
      memory_array[7052] <= 3'b000;
      memory_array[7053] <= 3'b000;
      memory_array[7054] <= 3'b101;
      memory_array[7055] <= 3'b000;
      memory_array[7056] <= 3'b000;
      memory_array[7057] <= 3'b000;
      memory_array[7058] <= 3'b101;
      memory_array[7059] <= 3'b000;
      memory_array[7060] <= 3'b101;
      memory_array[7061] <= 3'b101;
      memory_array[7062] <= 3'b101;
      memory_array[7063] <= 3'b000;
      memory_array[7064] <= 3'b101;
      memory_array[7065] <= 3'b101;
      memory_array[7066] <= 3'b101;
      memory_array[7067] <= 3'b101;
      memory_array[7068] <= 3'b101;
      memory_array[7069] <= 3'b101;
      memory_array[7070] <= 3'b101;
      memory_array[7071] <= 3'b101;
      memory_array[7072] <= 3'b101;
      memory_array[7073] <= 3'b000;
      memory_array[7074] <= 3'b101;
      memory_array[7075] <= 3'b000;
      memory_array[7076] <= 3'b101;
      memory_array[7077] <= 3'b101;
      memory_array[7078] <= 3'b000;
      memory_array[7079] <= 3'b101;
      memory_array[7080] <= 3'b101;
      memory_array[7081] <= 3'b101;
      memory_array[7082] <= 3'b000;
      memory_array[7083] <= 3'b000;
      memory_array[7084] <= 3'b101;
      memory_array[7085] <= 3'b000;
      memory_array[7086] <= 3'b111;
      memory_array[7087] <= 3'b111;
      memory_array[7088] <= 3'b111;
      memory_array[7089] <= 3'b000;
      memory_array[7090] <= 3'b000;
      memory_array[7091] <= 3'b101;
      memory_array[7092] <= 3'b111;
      memory_array[7093] <= 3'b111;
      memory_array[7094] <= 3'b111;
      memory_array[7095] <= 3'b111;
      memory_array[7096] <= 3'b101;
      memory_array[7097] <= 3'b101;
      memory_array[7098] <= 3'b000;
      memory_array[7099] <= 3'b101;
      memory_array[7100] <= 3'b000;
      memory_array[7101] <= 3'b101;
      memory_array[7102] <= 3'b000;
      memory_array[7103] <= 3'b000;
      memory_array[7104] <= 3'b101;
      memory_array[7105] <= 3'b000;
      memory_array[7106] <= 3'b101;
      memory_array[7107] <= 3'b101;
      memory_array[7108] <= 3'b000;
      memory_array[7109] <= 3'b101;
      memory_array[7110] <= 3'b101;
      memory_array[7111] <= 3'b000;
      memory_array[7112] <= 3'b000;
      memory_array[7113] <= 3'b000;
      memory_array[7114] <= 3'b000;
      memory_array[7115] <= 3'b101;
      memory_array[7116] <= 3'b000;
      memory_array[7117] <= 3'b101;
      memory_array[7118] <= 3'b101;
      memory_array[7119] <= 3'b101;
      memory_array[7120] <= 3'b101;
      memory_array[7121] <= 3'b000;
      memory_array[7122] <= 3'b101;
      memory_array[7123] <= 3'b101;
      memory_array[7124] <= 3'b000;
      memory_array[7125] <= 3'b101;
      memory_array[7126] <= 3'b000;
      memory_array[7127] <= 3'b101;
      memory_array[7128] <= 3'b101;
      memory_array[7129] <= 3'b101;
      memory_array[7130] <= 3'b101;
      memory_array[7131] <= 3'b101;
      memory_array[7132] <= 3'b101;
      memory_array[7133] <= 3'b101;
      memory_array[7134] <= 3'b101;
      memory_array[7135] <= 3'b101;
      memory_array[7136] <= 3'b000;
      memory_array[7137] <= 3'b000;
      memory_array[7138] <= 3'b101;
      memory_array[7139] <= 3'b101;
      memory_array[7140] <= 3'b000;
      memory_array[7141] <= 3'b101;
      memory_array[7142] <= 3'b101;
      memory_array[7143] <= 3'b000;
      memory_array[7144] <= 3'b000;
      memory_array[7145] <= 3'b101;
      memory_array[7146] <= 3'b000;
      memory_array[7147] <= 3'b000;
      memory_array[7148] <= 3'b000;
      memory_array[7149] <= 3'b101;
      memory_array[7150] <= 3'b000;
      memory_array[7151] <= 3'b000;
      memory_array[7152] <= 3'b101;
      memory_array[7153] <= 3'b111;
      memory_array[7154] <= 3'b111;
      memory_array[7155] <= 3'b111;
      memory_array[7156] <= 3'b111;
      memory_array[7157] <= 3'b101;
      memory_array[7158] <= 3'b000;
      memory_array[7159] <= 3'b000;
      memory_array[7160] <= 3'b111;
      memory_array[7161] <= 3'b000;
      memory_array[7162] <= 3'b101;
      memory_array[7163] <= 3'b000;
      memory_array[7164] <= 3'b110;
      memory_array[7165] <= 3'b000;
      memory_array[7166] <= 3'b101;
      memory_array[7167] <= 3'b000;
      memory_array[7168] <= 3'b110;
      memory_array[7169] <= 3'b000;
      memory_array[7170] <= 3'b101;
      memory_array[7171] <= 3'b000;
      memory_array[7172] <= 3'b000;
      memory_array[7173] <= 3'b110;
      memory_array[7174] <= 3'b110;
      memory_array[7175] <= 3'b000;
      memory_array[7176] <= 3'b000;
      memory_array[7177] <= 3'b101;
      memory_array[7178] <= 3'b000;
      memory_array[7179] <= 3'b110;
      memory_array[7180] <= 3'b000;
      memory_array[7181] <= 3'b000;
      memory_array[7182] <= 3'b000;
      memory_array[7183] <= 3'b110;
      memory_array[7184] <= 3'b101;
      memory_array[7185] <= 3'b101;
      memory_array[7186] <= 3'b000;
      memory_array[7187] <= 3'b101;
      memory_array[7188] <= 3'b000;
      memory_array[7189] <= 3'b000;
      memory_array[7190] <= 3'b000;
      memory_array[7191] <= 3'b101;
      memory_array[7192] <= 3'b101;
      memory_array[7193] <= 3'b101;
      memory_array[7194] <= 3'b101;
      memory_array[7195] <= 3'b101;
      memory_array[7196] <= 3'b101;
      memory_array[7197] <= 3'b101;
      memory_array[7198] <= 3'b101;
      memory_array[7199] <= 3'b101;
      memory_array[7200] <= 3'b000;
      memory_array[7201] <= 3'b000;
      memory_array[7202] <= 3'b000;
      memory_array[7203] <= 3'b110;
      memory_array[7204] <= 3'b110;
      memory_array[7205] <= 3'b000;
      memory_array[7206] <= 3'b000;
      memory_array[7207] <= 3'b000;
      memory_array[7208] <= 3'b101;
      memory_array[7209] <= 3'b000;
      memory_array[7210] <= 3'b000;
      memory_array[7211] <= 3'b000;
      memory_array[7212] <= 3'b000;
      memory_array[7213] <= 3'b000;
      memory_array[7214] <= 3'b110;
      memory_array[7215] <= 3'b000;
      memory_array[7216] <= 3'b000;
      memory_array[7217] <= 3'b000;
      memory_array[7218] <= 3'b110;
      memory_array[7219] <= 3'b000;
      memory_array[7220] <= 3'b101;
      memory_array[7221] <= 3'b000;
      memory_array[7222] <= 3'b000;
      memory_array[7223] <= 3'b110;
      memory_array[7224] <= 3'b000;
      memory_array[7225] <= 3'b101;
      memory_array[7226] <= 3'b000;
      memory_array[7227] <= 3'b101;
      memory_array[7228] <= 3'b000;
      memory_array[7229] <= 3'b000;
      memory_array[7230] <= 3'b101;
      memory_array[7231] <= 3'b101;
      memory_array[7232] <= 3'b000;
      memory_array[7233] <= 3'b000;
      memory_array[7234] <= 3'b110;
      memory_array[7235] <= 3'b000;
      memory_array[7236] <= 3'b000;
      memory_array[7237] <= 3'b000;
      memory_array[7238] <= 3'b101;
      memory_array[7239] <= 3'b101;
      memory_array[7240] <= 3'b000;
      memory_array[7241] <= 3'b111;
      memory_array[7242] <= 3'b111;
      memory_array[7243] <= 3'b111;
      memory_array[7244] <= 3'b111;
      memory_array[7245] <= 3'b111;
      memory_array[7246] <= 3'b000;
      memory_array[7247] <= 3'b101;
      memory_array[7248] <= 3'b000;
      memory_array[7249] <= 3'b000;
      memory_array[7250] <= 3'b000;
      memory_array[7251] <= 3'b000;
      memory_array[7252] <= 3'b101;
      memory_array[7253] <= 3'b101;
      memory_array[7254] <= 3'b000;
      memory_array[7255] <= 3'b101;
      memory_array[7256] <= 3'b101;
      memory_array[7257] <= 3'b101;
      memory_array[7258] <= 3'b000;
      memory_array[7259] <= 3'b101;
      memory_array[7260] <= 3'b000;
      memory_array[7261] <= 3'b101;
      memory_array[7262] <= 3'b101;
      memory_array[7263] <= 3'b101;
      memory_array[7264] <= 3'b101;
      memory_array[7265] <= 3'b101;
      memory_array[7266] <= 3'b000;
      memory_array[7267] <= 3'b101;
      memory_array[7268] <= 3'b101;
      memory_array[7269] <= 3'b101;
      memory_array[7270] <= 3'b101;
      memory_array[7271] <= 3'b101;
      memory_array[7272] <= 3'b101;
      memory_array[7273] <= 3'b101;
      memory_array[7274] <= 3'b000;
      memory_array[7275] <= 3'b101;
      memory_array[7276] <= 3'b101;
      memory_array[7277] <= 3'b000;
      memory_array[7278] <= 3'b101;
      memory_array[7279] <= 3'b000;
      memory_array[7280] <= 3'b101;
      memory_array[7281] <= 3'b101;
      memory_array[7282] <= 3'b000;
      memory_array[7283] <= 3'b101;
      memory_array[7284] <= 3'b000;
      memory_array[7285] <= 3'b101;
      memory_array[7286] <= 3'b111;
      memory_array[7287] <= 3'b111;
      memory_array[7288] <= 3'b111;
      memory_array[7289] <= 3'b000;
      memory_array[7290] <= 3'b000;
      memory_array[7291] <= 3'b101;
      memory_array[7292] <= 3'b111;
      memory_array[7293] <= 3'b111;
      memory_array[7294] <= 3'b111;
      memory_array[7295] <= 3'b111;
      memory_array[7296] <= 3'b000;
      memory_array[7297] <= 3'b111;
      memory_array[7298] <= 3'b000;
      memory_array[7299] <= 3'b101;
      memory_array[7300] <= 3'b101;
      memory_array[7301] <= 3'b111;
      memory_array[7302] <= 3'b101;
      memory_array[7303] <= 3'b000;
      memory_array[7304] <= 3'b101;
      memory_array[7305] <= 3'b101;
      memory_array[7306] <= 3'b101;
      memory_array[7307] <= 3'b101;
      memory_array[7308] <= 3'b101;
      memory_array[7309] <= 3'b000;
      memory_array[7310] <= 3'b101;
      memory_array[7311] <= 3'b101;
      memory_array[7312] <= 3'b000;
      memory_array[7313] <= 3'b101;
      memory_array[7314] <= 3'b101;
      memory_array[7315] <= 3'b000;
      memory_array[7316] <= 3'b101;
      memory_array[7317] <= 3'b000;
      memory_array[7318] <= 3'b101;
      memory_array[7319] <= 3'b101;
      memory_array[7320] <= 3'b000;
      memory_array[7321] <= 3'b101;
      memory_array[7322] <= 3'b000;
      memory_array[7323] <= 3'b101;
      memory_array[7324] <= 3'b101;
      memory_array[7325] <= 3'b000;
      memory_array[7326] <= 3'b101;
      memory_array[7327] <= 3'b101;
      memory_array[7328] <= 3'b101;
      memory_array[7329] <= 3'b101;
      memory_array[7330] <= 3'b101;
      memory_array[7331] <= 3'b101;
      memory_array[7332] <= 3'b000;
      memory_array[7333] <= 3'b000;
      memory_array[7334] <= 3'b101;
      memory_array[7335] <= 3'b101;
      memory_array[7336] <= 3'b101;
      memory_array[7337] <= 3'b000;
      memory_array[7338] <= 3'b101;
      memory_array[7339] <= 3'b000;
      memory_array[7340] <= 3'b101;
      memory_array[7341] <= 3'b000;
      memory_array[7342] <= 3'b101;
      memory_array[7343] <= 3'b101;
      memory_array[7344] <= 3'b101;
      memory_array[7345] <= 3'b000;
      memory_array[7346] <= 3'b101;
      memory_array[7347] <= 3'b101;
      memory_array[7348] <= 3'b000;
      memory_array[7349] <= 3'b000;
      memory_array[7350] <= 3'b000;
      memory_array[7351] <= 3'b000;
      memory_array[7352] <= 3'b000;
      memory_array[7353] <= 3'b000;
      memory_array[7354] <= 3'b111;
      memory_array[7355] <= 3'b111;
      memory_array[7356] <= 3'b111;
      memory_array[7357] <= 3'b111;
      memory_array[7358] <= 3'b111;
      memory_array[7359] <= 3'b000;
      memory_array[7360] <= 3'b101;
      memory_array[7361] <= 3'b101;
      memory_array[7362] <= 3'b101;
      memory_array[7363] <= 3'b000;
      memory_array[7364] <= 3'b000;
      memory_array[7365] <= 3'b000;
      memory_array[7366] <= 3'b000;
      memory_array[7367] <= 3'b000;
      memory_array[7368] <= 3'b101;
      memory_array[7369] <= 3'b101;
      memory_array[7370] <= 3'b000;
      memory_array[7371] <= 3'b000;
      memory_array[7372] <= 3'b101;
      memory_array[7373] <= 3'b000;
      memory_array[7374] <= 3'b101;
      memory_array[7375] <= 3'b000;
      memory_array[7376] <= 3'b000;
      memory_array[7377] <= 3'b000;
      memory_array[7378] <= 3'b000;
      memory_array[7379] <= 3'b101;
      memory_array[7380] <= 3'b000;
      memory_array[7381] <= 3'b000;
      memory_array[7382] <= 3'b000;
      memory_array[7383] <= 3'b110;
      memory_array[7384] <= 3'b110;
      memory_array[7385] <= 3'b000;
      memory_array[7386] <= 3'b000;
      memory_array[7387] <= 3'b000;
      memory_array[7388] <= 3'b000;
      memory_array[7389] <= 3'b000;
      memory_array[7390] <= 3'b000;
      memory_array[7391] <= 3'b101;
      memory_array[7392] <= 3'b000;
      memory_array[7393] <= 3'b110;
      memory_array[7394] <= 3'b110;
      memory_array[7395] <= 3'b000;
      memory_array[7396] <= 3'b000;
      memory_array[7397] <= 3'b000;
      memory_array[7398] <= 3'b110;
      memory_array[7399] <= 3'b110;
      memory_array[7400] <= 3'b101;
      memory_array[7401] <= 3'b000;
      memory_array[7402] <= 3'b000;
      memory_array[7403] <= 3'b110;
      memory_array[7404] <= 3'b110;
      memory_array[7405] <= 3'b000;
      memory_array[7406] <= 3'b000;
      memory_array[7407] <= 3'b101;
      memory_array[7408] <= 3'b101;
      memory_array[7409] <= 3'b000;
      memory_array[7410] <= 3'b000;
      memory_array[7411] <= 3'b000;
      memory_array[7412] <= 3'b101;
      memory_array[7413] <= 3'b000;
      memory_array[7414] <= 3'b101;
      memory_array[7415] <= 3'b111;
      memory_array[7416] <= 3'b000;
      memory_array[7417] <= 3'b000;
      memory_array[7418] <= 3'b000;
      memory_array[7419] <= 3'b000;
      memory_array[7420] <= 3'b000;
      memory_array[7421] <= 3'b000;
      memory_array[7422] <= 3'b000;
      memory_array[7423] <= 3'b110;
      memory_array[7424] <= 3'b101;
      memory_array[7425] <= 3'b101;
      memory_array[7426] <= 3'b000;
      memory_array[7427] <= 3'b000;
      memory_array[7428] <= 3'b110;
      memory_array[7429] <= 3'b000;
      memory_array[7430] <= 3'b101;
      memory_array[7431] <= 3'b000;
      memory_array[7432] <= 3'b000;
      memory_array[7433] <= 3'b000;
      memory_array[7434] <= 3'b000;
      memory_array[7435] <= 3'b000;
      memory_array[7436] <= 3'b000;
      memory_array[7437] <= 3'b000;
      memory_array[7438] <= 3'b101;
      memory_array[7439] <= 3'b101;
      memory_array[7440] <= 3'b111;
      memory_array[7441] <= 3'b111;
      memory_array[7442] <= 3'b111;
      memory_array[7443] <= 3'b111;
      memory_array[7444] <= 3'b101;
      memory_array[7445] <= 3'b000;
      memory_array[7446] <= 3'b101;
      memory_array[7447] <= 3'b101;
      memory_array[7448] <= 3'b101;
      memory_array[7449] <= 3'b000;
      memory_array[7450] <= 3'b000;
      memory_array[7451] <= 3'b000;
      memory_array[7452] <= 3'b000;
      memory_array[7453] <= 3'b101;
      memory_array[7454] <= 3'b101;
      memory_array[7455] <= 3'b000;
      memory_array[7456] <= 3'b000;
      memory_array[7457] <= 3'b000;
      memory_array[7458] <= 3'b101;
      memory_array[7459] <= 3'b000;
      memory_array[7460] <= 3'b101;
      memory_array[7461] <= 3'b101;
      memory_array[7462] <= 3'b000;
      memory_array[7463] <= 3'b101;
      memory_array[7464] <= 3'b101;
      memory_array[7465] <= 3'b101;
      memory_array[7466] <= 3'b101;
      memory_array[7467] <= 3'b000;
      memory_array[7468] <= 3'b101;
      memory_array[7469] <= 3'b101;
      memory_array[7470] <= 3'b101;
      memory_array[7471] <= 3'b101;
      memory_array[7472] <= 3'b101;
      memory_array[7473] <= 3'b101;
      memory_array[7474] <= 3'b000;
      memory_array[7475] <= 3'b000;
      memory_array[7476] <= 3'b101;
      memory_array[7477] <= 3'b101;
      memory_array[7478] <= 3'b000;
      memory_array[7479] <= 3'b101;
      memory_array[7480] <= 3'b101;
      memory_array[7481] <= 3'b101;
      memory_array[7482] <= 3'b000;
      memory_array[7483] <= 3'b101;
      memory_array[7484] <= 3'b101;
      memory_array[7485] <= 3'b111;
      memory_array[7486] <= 3'b101;
      memory_array[7487] <= 3'b111;
      memory_array[7488] <= 3'b000;
      memory_array[7489] <= 3'b101;
      memory_array[7490] <= 3'b101;
      memory_array[7491] <= 3'b101;
      memory_array[7492] <= 3'b101;
      memory_array[7493] <= 3'b111;
      memory_array[7494] <= 3'b000;
      memory_array[7495] <= 3'b101;
      memory_array[7496] <= 3'b101;
      memory_array[7497] <= 3'b111;
      memory_array[7498] <= 3'b111;
      memory_array[7499] <= 3'b000;
      memory_array[7500] <= 3'b101;
      memory_array[7501] <= 3'b111;
      memory_array[7502] <= 3'b111;
      memory_array[7503] <= 3'b101;
      memory_array[7504] <= 3'b101;
      memory_array[7505] <= 3'b000;
      memory_array[7506] <= 3'b000;
      memory_array[7507] <= 3'b101;
      memory_array[7508] <= 3'b101;
      memory_array[7509] <= 3'b101;
      memory_array[7510] <= 3'b101;
      memory_array[7511] <= 3'b101;
      memory_array[7512] <= 3'b101;
      memory_array[7513] <= 3'b101;
      memory_array[7514] <= 3'b101;
      memory_array[7515] <= 3'b101;
      memory_array[7516] <= 3'b101;
      memory_array[7517] <= 3'b000;
      memory_array[7518] <= 3'b101;
      memory_array[7519] <= 3'b101;
      memory_array[7520] <= 3'b101;
      memory_array[7521] <= 3'b000;
      memory_array[7522] <= 3'b000;
      memory_array[7523] <= 3'b101;
      memory_array[7524] <= 3'b000;
      memory_array[7525] <= 3'b000;
      memory_array[7526] <= 3'b101;
      memory_array[7527] <= 3'b101;
      memory_array[7528] <= 3'b101;
      memory_array[7529] <= 3'b101;
      memory_array[7530] <= 3'b101;
      memory_array[7531] <= 3'b101;
      memory_array[7532] <= 3'b101;
      memory_array[7533] <= 3'b101;
      memory_array[7534] <= 3'b101;
      memory_array[7535] <= 3'b101;
      memory_array[7536] <= 3'b101;
      memory_array[7537] <= 3'b101;
      memory_array[7538] <= 3'b101;
      memory_array[7539] <= 3'b101;
      memory_array[7540] <= 3'b000;
      memory_array[7541] <= 3'b101;
      memory_array[7542] <= 3'b000;
      memory_array[7543] <= 3'b000;
      memory_array[7544] <= 3'b000;
      memory_array[7545] <= 3'b101;
      memory_array[7546] <= 3'b101;
      memory_array[7547] <= 3'b101;
      memory_array[7548] <= 3'b000;
      memory_array[7549] <= 3'b000;
      memory_array[7550] <= 3'b000;
      memory_array[7551] <= 3'b101;
      memory_array[7552] <= 3'b101;
      memory_array[7553] <= 3'b101;
      memory_array[7554] <= 3'b000;
      memory_array[7555] <= 3'b101;
      memory_array[7556] <= 3'b111;
      memory_array[7557] <= 3'b111;
      memory_array[7558] <= 3'b111;
      memory_array[7559] <= 3'b111;
      memory_array[7560] <= 3'b101;
      memory_array[7561] <= 3'b101;
      memory_array[7562] <= 3'b101;
      memory_array[7563] <= 3'b000;
      memory_array[7564] <= 3'b110;
      memory_array[7565] <= 3'b000;
      memory_array[7566] <= 3'b000;
      memory_array[7567] <= 3'b000;
      memory_array[7568] <= 3'b000;
      memory_array[7569] <= 3'b101;
      memory_array[7570] <= 3'b000;
      memory_array[7571] <= 3'b000;
      memory_array[7572] <= 3'b101;
      memory_array[7573] <= 3'b000;
      memory_array[7574] <= 3'b101;
      memory_array[7575] <= 3'b101;
      memory_array[7576] <= 3'b000;
      memory_array[7577] <= 3'b000;
      memory_array[7578] <= 3'b110;
      memory_array[7579] <= 3'b110;
      memory_array[7580] <= 3'b000;
      memory_array[7581] <= 3'b000;
      memory_array[7582] <= 3'b000;
      memory_array[7583] <= 3'b000;
      memory_array[7584] <= 3'b111;
      memory_array[7585] <= 3'b101;
      memory_array[7586] <= 3'b000;
      memory_array[7587] <= 3'b101;
      memory_array[7588] <= 3'b000;
      memory_array[7589] <= 3'b000;
      memory_array[7590] <= 3'b000;
      memory_array[7591] <= 3'b101;
      memory_array[7592] <= 3'b101;
      memory_array[7593] <= 3'b110;
      memory_array[7594] <= 3'b110;
      memory_array[7595] <= 3'b000;
      memory_array[7596] <= 3'b000;
      memory_array[7597] <= 3'b000;
      memory_array[7598] <= 3'b110;
      memory_array[7599] <= 3'b101;
      memory_array[7600] <= 3'b101;
      memory_array[7601] <= 3'b101;
      memory_array[7602] <= 3'b110;
      memory_array[7603] <= 3'b101;
      memory_array[7604] <= 3'b101;
      memory_array[7605] <= 3'b110;
      memory_array[7606] <= 3'b101;
      memory_array[7607] <= 3'b101;
      memory_array[7608] <= 3'b101;
      memory_array[7609] <= 3'b000;
      memory_array[7610] <= 3'b000;
      memory_array[7611] <= 3'b101;
      memory_array[7612] <= 3'b000;
      memory_array[7613] <= 3'b000;
      memory_array[7614] <= 3'b000;
      memory_array[7615] <= 3'b101;
      memory_array[7616] <= 3'b110;
      memory_array[7617] <= 3'b110;
      memory_array[7618] <= 3'b000;
      memory_array[7619] <= 3'b000;
      memory_array[7620] <= 3'b110;
      memory_array[7621] <= 3'b110;
      memory_array[7622] <= 3'b110;
      memory_array[7623] <= 3'b000;
      memory_array[7624] <= 3'b101;
      memory_array[7625] <= 3'b101;
      memory_array[7626] <= 3'b000;
      memory_array[7627] <= 3'b110;
      memory_array[7628] <= 3'b000;
      memory_array[7629] <= 3'b000;
      memory_array[7630] <= 3'b000;
      memory_array[7631] <= 3'b110;
      memory_array[7632] <= 3'b110;
      memory_array[7633] <= 3'b000;
      memory_array[7634] <= 3'b000;
      memory_array[7635] <= 3'b000;
      memory_array[7636] <= 3'b101;
      memory_array[7637] <= 3'b101;
      memory_array[7638] <= 3'b000;
      memory_array[7639] <= 3'b111;
      memory_array[7640] <= 3'b111;
      memory_array[7641] <= 3'b111;
      memory_array[7642] <= 3'b111;
      memory_array[7643] <= 3'b111;
      memory_array[7644] <= 3'b000;
      memory_array[7645] <= 3'b101;
      memory_array[7646] <= 3'b101;
      memory_array[7647] <= 3'b101;
      memory_array[7648] <= 3'b101;
      memory_array[7649] <= 3'b101;
      memory_array[7650] <= 3'b000;
      memory_array[7651] <= 3'b101;
      memory_array[7652] <= 3'b101;
      memory_array[7653] <= 3'b101;
      memory_array[7654] <= 3'b101;
      memory_array[7655] <= 3'b000;
      memory_array[7656] <= 3'b000;
      memory_array[7657] <= 3'b101;
      memory_array[7658] <= 3'b000;
      memory_array[7659] <= 3'b101;
      memory_array[7660] <= 3'b101;
      memory_array[7661] <= 3'b101;
      memory_array[7662] <= 3'b101;
      memory_array[7663] <= 3'b101;
      memory_array[7664] <= 3'b101;
      memory_array[7665] <= 3'b000;
      memory_array[7666] <= 3'b101;
      memory_array[7667] <= 3'b101;
      memory_array[7668] <= 3'b000;
      memory_array[7669] <= 3'b101;
      memory_array[7670] <= 3'b101;
      memory_array[7671] <= 3'b101;
      memory_array[7672] <= 3'b101;
      memory_array[7673] <= 3'b000;
      memory_array[7674] <= 3'b101;
      memory_array[7675] <= 3'b101;
      memory_array[7676] <= 3'b101;
      memory_array[7677] <= 3'b101;
      memory_array[7678] <= 3'b000;
      memory_array[7679] <= 3'b101;
      memory_array[7680] <= 3'b101;
      memory_array[7681] <= 3'b101;
      memory_array[7682] <= 3'b101;
      memory_array[7683] <= 3'b101;
      memory_array[7684] <= 3'b101;
      memory_array[7685] <= 3'b111;
      memory_array[7686] <= 3'b101;
      memory_array[7687] <= 3'b111;
      memory_array[7688] <= 3'b000;
      memory_array[7689] <= 3'b101;
      memory_array[7690] <= 3'b101;
      memory_array[7691] <= 3'b101;
      memory_array[7692] <= 3'b000;
      memory_array[7693] <= 3'b111;
      memory_array[7694] <= 3'b000;
      memory_array[7695] <= 3'b101;
      memory_array[7696] <= 3'b101;
      memory_array[7697] <= 3'b000;
      memory_array[7698] <= 3'b111;
      memory_array[7699] <= 3'b101;
      memory_array[7700] <= 3'b101;
      memory_array[7701] <= 3'b111;
      memory_array[7702] <= 3'b101;
      memory_array[7703] <= 3'b000;
      memory_array[7704] <= 3'b101;
      memory_array[7705] <= 3'b101;
      memory_array[7706] <= 3'b101;
      memory_array[7707] <= 3'b000;
      memory_array[7708] <= 3'b101;
      memory_array[7709] <= 3'b101;
      memory_array[7710] <= 3'b000;
      memory_array[7711] <= 3'b101;
      memory_array[7712] <= 3'b000;
      memory_array[7713] <= 3'b101;
      memory_array[7714] <= 3'b101;
      memory_array[7715] <= 3'b101;
      memory_array[7716] <= 3'b101;
      memory_array[7717] <= 3'b101;
      memory_array[7718] <= 3'b101;
      memory_array[7719] <= 3'b101;
      memory_array[7720] <= 3'b101;
      memory_array[7721] <= 3'b000;
      memory_array[7722] <= 3'b101;
      memory_array[7723] <= 3'b101;
      memory_array[7724] <= 3'b101;
      memory_array[7725] <= 3'b101;
      memory_array[7726] <= 3'b000;
      memory_array[7727] <= 3'b101;
      memory_array[7728] <= 3'b101;
      memory_array[7729] <= 3'b101;
      memory_array[7730] <= 3'b101;
      memory_array[7731] <= 3'b000;
      memory_array[7732] <= 3'b101;
      memory_array[7733] <= 3'b101;
      memory_array[7734] <= 3'b000;
      memory_array[7735] <= 3'b101;
      memory_array[7736] <= 3'b101;
      memory_array[7737] <= 3'b000;
      memory_array[7738] <= 3'b101;
      memory_array[7739] <= 3'b101;
      memory_array[7740] <= 3'b101;
      memory_array[7741] <= 3'b000;
      memory_array[7742] <= 3'b101;
      memory_array[7743] <= 3'b000;
      memory_array[7744] <= 3'b000;
      memory_array[7745] <= 3'b101;
      memory_array[7746] <= 3'b101;
      memory_array[7747] <= 3'b101;
      memory_array[7748] <= 3'b101;
      memory_array[7749] <= 3'b000;
      memory_array[7750] <= 3'b101;
      memory_array[7751] <= 3'b101;
      memory_array[7752] <= 3'b000;
      memory_array[7753] <= 3'b101;
      memory_array[7754] <= 3'b000;
      memory_array[7755] <= 3'b000;
      memory_array[7756] <= 3'b111;
      memory_array[7757] <= 3'b111;
      memory_array[7758] <= 3'b111;
      memory_array[7759] <= 3'b111;
      memory_array[7760] <= 3'b111;
      memory_array[7761] <= 3'b000;
      memory_array[7762] <= 3'b000;
      memory_array[7763] <= 3'b101;
      memory_array[7764] <= 3'b000;
      memory_array[7765] <= 3'b110;
      memory_array[7766] <= 3'b110;
      memory_array[7767] <= 3'b110;
      memory_array[7768] <= 3'b000;
      memory_array[7769] <= 3'b000;
      memory_array[7770] <= 3'b000;
      memory_array[7771] <= 3'b110;
      memory_array[7772] <= 3'b110;
      memory_array[7773] <= 3'b000;
      memory_array[7774] <= 3'b101;
      memory_array[7775] <= 3'b101;
      memory_array[7776] <= 3'b110;
      memory_array[7777] <= 3'b110;
      memory_array[7778] <= 3'b000;
      memory_array[7779] <= 3'b000;
      memory_array[7780] <= 3'b110;
      memory_array[7781] <= 3'b110;
      memory_array[7782] <= 3'b110;
      memory_array[7783] <= 3'b000;
      memory_array[7784] <= 3'b101;
      memory_array[7785] <= 3'b000;
      memory_array[7786] <= 3'b000;
      memory_array[7787] <= 3'b101;
      memory_array[7788] <= 3'b101;
      memory_array[7789] <= 3'b000;
      memory_array[7790] <= 3'b000;
      memory_array[7791] <= 3'b101;
      memory_array[7792] <= 3'b101;
      memory_array[7793] <= 3'b101;
      memory_array[7794] <= 3'b000;
      memory_array[7795] <= 3'b101;
      memory_array[7796] <= 3'b101;
      memory_array[7797] <= 3'b110;
      memory_array[7798] <= 3'b101;
      memory_array[7799] <= 3'b101;
      memory_array[7800] <= 3'b101;
      memory_array[7801] <= 3'b101;
      memory_array[7802] <= 3'b101;
      memory_array[7803] <= 3'b111;
      memory_array[7804] <= 3'b111;
      memory_array[7805] <= 3'b101;
      memory_array[7806] <= 3'b101;
      memory_array[7807] <= 3'b101;
      memory_array[7808] <= 3'b101;
      memory_array[7809] <= 3'b000;
      memory_array[7810] <= 3'b000;
      memory_array[7811] <= 3'b000;
      memory_array[7812] <= 3'b000;
      memory_array[7813] <= 3'b110;
      memory_array[7814] <= 3'b000;
      memory_array[7815] <= 3'b000;
      memory_array[7816] <= 3'b000;
      memory_array[7817] <= 3'b000;
      memory_array[7818] <= 3'b110;
      memory_array[7819] <= 3'b110;
      memory_array[7820] <= 3'b000;
      memory_array[7821] <= 3'b000;
      memory_array[7822] <= 3'b000;
      memory_array[7823] <= 3'b110;
      memory_array[7824] <= 3'b000;
      memory_array[7825] <= 3'b101;
      memory_array[7826] <= 3'b000;
      memory_array[7827] <= 3'b000;
      memory_array[7828] <= 3'b110;
      memory_array[7829] <= 3'b000;
      memory_array[7830] <= 3'b000;
      memory_array[7831] <= 3'b000;
      memory_array[7832] <= 3'b000;
      memory_array[7833] <= 3'b110;
      memory_array[7834] <= 3'b110;
      memory_array[7835] <= 3'b000;
      memory_array[7836] <= 3'b000;
      memory_array[7837] <= 3'b000;
      memory_array[7838] <= 3'b101;
      memory_array[7839] <= 3'b111;
      memory_array[7840] <= 3'b111;
      memory_array[7841] <= 3'b111;
      memory_array[7842] <= 3'b111;
      memory_array[7843] <= 3'b101;
      memory_array[7844] <= 3'b101;
      memory_array[7845] <= 3'b101;
      memory_array[7846] <= 3'b000;
      memory_array[7847] <= 3'b101;
      memory_array[7848] <= 3'b101;
      memory_array[7849] <= 3'b101;
      memory_array[7850] <= 3'b101;
      memory_array[7851] <= 3'b101;
      memory_array[7852] <= 3'b101;
      memory_array[7853] <= 3'b000;
      memory_array[7854] <= 3'b101;
      memory_array[7855] <= 3'b000;
      memory_array[7856] <= 3'b111;
      memory_array[7857] <= 3'b101;
      memory_array[7858] <= 3'b000;
      memory_array[7859] <= 3'b000;
      memory_array[7860] <= 3'b000;
      memory_array[7861] <= 3'b000;
      memory_array[7862] <= 3'b101;
      memory_array[7863] <= 3'b101;
      memory_array[7864] <= 3'b101;
      memory_array[7865] <= 3'b101;
      memory_array[7866] <= 3'b101;
      memory_array[7867] <= 3'b101;
      memory_array[7868] <= 3'b101;
      memory_array[7869] <= 3'b101;
      memory_array[7870] <= 3'b101;
      memory_array[7871] <= 3'b101;
      memory_array[7872] <= 3'b101;
      memory_array[7873] <= 3'b000;
      memory_array[7874] <= 3'b101;
      memory_array[7875] <= 3'b101;
      memory_array[7876] <= 3'b101;
      memory_array[7877] <= 3'b101;
      memory_array[7878] <= 3'b101;
      memory_array[7879] <= 3'b101;
      memory_array[7880] <= 3'b101;
      memory_array[7881] <= 3'b101;
      memory_array[7882] <= 3'b101;
      memory_array[7883] <= 3'b101;
      memory_array[7884] <= 3'b111;
      memory_array[7885] <= 3'b111;
      memory_array[7886] <= 3'b101;
      memory_array[7887] <= 3'b101;
      memory_array[7888] <= 3'b101;
      memory_array[7889] <= 3'b101;
      memory_array[7890] <= 3'b000;
      memory_array[7891] <= 3'b000;
      memory_array[7892] <= 3'b101;
      memory_array[7893] <= 3'b111;
      memory_array[7894] <= 3'b000;
      memory_array[7895] <= 3'b000;
      memory_array[7896] <= 3'b101;
      memory_array[7897] <= 3'b000;
      memory_array[7898] <= 3'b111;
      memory_array[7899] <= 3'b101;
      memory_array[7900] <= 3'b101;
      memory_array[7901] <= 3'b000;
      memory_array[7902] <= 3'b000;
      memory_array[7903] <= 3'b101;
      memory_array[7904] <= 3'b101;
      memory_array[7905] <= 3'b000;
      memory_array[7906] <= 3'b101;
      memory_array[7907] <= 3'b000;
      memory_array[7908] <= 3'b000;
      memory_array[7909] <= 3'b101;
      memory_array[7910] <= 3'b101;
      memory_array[7911] <= 3'b101;
      memory_array[7912] <= 3'b101;
      memory_array[7913] <= 3'b101;
      memory_array[7914] <= 3'b101;
      memory_array[7915] <= 3'b101;
      memory_array[7916] <= 3'b101;
      memory_array[7917] <= 3'b000;
      memory_array[7918] <= 3'b101;
      memory_array[7919] <= 3'b101;
      memory_array[7920] <= 3'b101;
      memory_array[7921] <= 3'b101;
      memory_array[7922] <= 3'b101;
      memory_array[7923] <= 3'b101;
      memory_array[7924] <= 3'b101;
      memory_array[7925] <= 3'b101;
      memory_array[7926] <= 3'b000;
      memory_array[7927] <= 3'b000;
      memory_array[7928] <= 3'b101;
      memory_array[7929] <= 3'b101;
      memory_array[7930] <= 3'b101;
      memory_array[7931] <= 3'b101;
      memory_array[7932] <= 3'b000;
      memory_array[7933] <= 3'b101;
      memory_array[7934] <= 3'b101;
      memory_array[7935] <= 3'b101;
      memory_array[7936] <= 3'b101;
      memory_array[7937] <= 3'b000;
      memory_array[7938] <= 3'b000;
      memory_array[7939] <= 3'b000;
      memory_array[7940] <= 3'b000;
      memory_array[7941] <= 3'b000;
      memory_array[7942] <= 3'b101;
      memory_array[7943] <= 3'b000;
      memory_array[7944] <= 3'b000;
      memory_array[7945] <= 3'b101;
      memory_array[7946] <= 3'b000;
      memory_array[7947] <= 3'b101;
      memory_array[7948] <= 3'b101;
      memory_array[7949] <= 3'b101;
      memory_array[7950] <= 3'b101;
      memory_array[7951] <= 3'b101;
      memory_array[7952] <= 3'b000;
      memory_array[7953] <= 3'b000;
      memory_array[7954] <= 3'b101;
      memory_array[7955] <= 3'b000;
      memory_array[7956] <= 3'b101;
      memory_array[7957] <= 3'b111;
      memory_array[7958] <= 3'b111;
      memory_array[7959] <= 3'b111;
      memory_array[7960] <= 3'b111;
      memory_array[7961] <= 3'b101;
      memory_array[7962] <= 3'b101;
      memory_array[7963] <= 3'b000;
      memory_array[7964] <= 3'b000;
      memory_array[7965] <= 3'b000;
      memory_array[7966] <= 3'b000;
      memory_array[7967] <= 3'b000;
      memory_array[7968] <= 3'b110;
      memory_array[7969] <= 3'b000;
      memory_array[7970] <= 3'b000;
      memory_array[7971] <= 3'b000;
      memory_array[7972] <= 3'b000;
      memory_array[7973] <= 3'b000;
      memory_array[7974] <= 3'b101;
      memory_array[7975] <= 3'b000;
      memory_array[7976] <= 3'b000;
      memory_array[7977] <= 3'b000;
      memory_array[7978] <= 3'b110;
      memory_array[7979] <= 3'b110;
      memory_array[7980] <= 3'b000;
      memory_array[7981] <= 3'b000;
      memory_array[7982] <= 3'b000;
      memory_array[7983] <= 3'b110;
      memory_array[7984] <= 3'b110;
      memory_array[7985] <= 3'b000;
      memory_array[7986] <= 3'b000;
      memory_array[7987] <= 3'b000;
      memory_array[7988] <= 3'b000;
      memory_array[7989] <= 3'b000;
      memory_array[7990] <= 3'b000;
      memory_array[7991] <= 3'b101;
      memory_array[7992] <= 3'b101;
      memory_array[7993] <= 3'b101;
      memory_array[7994] <= 3'b101;
      memory_array[7995] <= 3'b111;
      memory_array[7996] <= 3'b111;
      memory_array[7997] <= 3'b101;
      memory_array[7998] <= 3'b101;
      memory_array[7999] <= 3'b101;
      memory_array[8000] <= 3'b101;
      memory_array[8001] <= 3'b101;
      memory_array[8002] <= 3'b101;
      memory_array[8003] <= 3'b101;
      memory_array[8004] <= 3'b101;
      memory_array[8005] <= 3'b101;
      memory_array[8006] <= 3'b101;
      memory_array[8007] <= 3'b101;
      memory_array[8008] <= 3'b101;
      memory_array[8009] <= 3'b000;
      memory_array[8010] <= 3'b000;
      memory_array[8011] <= 3'b110;
      memory_array[8012] <= 3'b000;
      memory_array[8013] <= 3'b101;
      memory_array[8014] <= 3'b000;
      memory_array[8015] <= 3'b110;
      memory_array[8016] <= 3'b110;
      memory_array[8017] <= 3'b110;
      memory_array[8018] <= 3'b000;
      memory_array[8019] <= 3'b000;
      memory_array[8020] <= 3'b110;
      memory_array[8021] <= 3'b110;
      memory_array[8022] <= 3'b110;
      memory_array[8023] <= 3'b000;
      memory_array[8024] <= 3'b000;
      memory_array[8025] <= 3'b000;
      memory_array[8026] <= 3'b101;
      memory_array[8027] <= 3'b110;
      memory_array[8028] <= 3'b000;
      memory_array[8029] <= 3'b000;
      memory_array[8030] <= 3'b110;
      memory_array[8031] <= 3'b110;
      memory_array[8032] <= 3'b110;
      memory_array[8033] <= 3'b000;
      memory_array[8034] <= 3'b000;
      memory_array[8035] <= 3'b110;
      memory_array[8036] <= 3'b000;
      memory_array[8037] <= 3'b101;
      memory_array[8038] <= 3'b111;
      memory_array[8039] <= 3'b111;
      memory_array[8040] <= 3'b111;
      memory_array[8041] <= 3'b111;
      memory_array[8042] <= 3'b101;
      memory_array[8043] <= 3'b000;
      memory_array[8044] <= 3'b101;
      memory_array[8045] <= 3'b101;
      memory_array[8046] <= 3'b000;
      memory_array[8047] <= 3'b000;
      memory_array[8048] <= 3'b101;
      memory_array[8049] <= 3'b101;
      memory_array[8050] <= 3'b000;
      memory_array[8051] <= 3'b101;
      memory_array[8052] <= 3'b101;
      memory_array[8053] <= 3'b101;
      memory_array[8054] <= 3'b101;
      memory_array[8055] <= 3'b101;
      memory_array[8056] <= 3'b111;
      memory_array[8057] <= 3'b101;
      memory_array[8058] <= 3'b101;
      memory_array[8059] <= 3'b101;
      memory_array[8060] <= 3'b000;
      memory_array[8061] <= 3'b101;
      memory_array[8062] <= 3'b101;
      memory_array[8063] <= 3'b101;
      memory_array[8064] <= 3'b101;
      memory_array[8065] <= 3'b101;
      memory_array[8066] <= 3'b101;
      memory_array[8067] <= 3'b101;
      memory_array[8068] <= 3'b101;
      memory_array[8069] <= 3'b101;
      memory_array[8070] <= 3'b101;
      memory_array[8071] <= 3'b000;
      memory_array[8072] <= 3'b000;
      memory_array[8073] <= 3'b101;
      memory_array[8074] <= 3'b101;
      memory_array[8075] <= 3'b101;
      memory_array[8076] <= 3'b000;
      memory_array[8077] <= 3'b000;
      memory_array[8078] <= 3'b101;
      memory_array[8079] <= 3'b000;
      memory_array[8080] <= 3'b101;
      memory_array[8081] <= 3'b101;
      memory_array[8082] <= 3'b000;
      memory_array[8083] <= 3'b111;
      memory_array[8084] <= 3'b111;
      memory_array[8085] <= 3'b111;
      memory_array[8086] <= 3'b111;
      memory_array[8087] <= 3'b101;
      memory_array[8088] <= 3'b000;
      memory_array[8089] <= 3'b000;
      memory_array[8090] <= 3'b000;
      memory_array[8091] <= 3'b111;
      memory_array[8092] <= 3'b101;
      memory_array[8093] <= 3'b111;
      memory_array[8094] <= 3'b000;
      memory_array[8095] <= 3'b101;
      memory_array[8096] <= 3'b101;
      memory_array[8097] <= 3'b111;
      memory_array[8098] <= 3'b111;
      memory_array[8099] <= 3'b000;
      memory_array[8100] <= 3'b000;
      memory_array[8101] <= 3'b101;
      memory_array[8102] <= 3'b000;
      memory_array[8103] <= 3'b000;
      memory_array[8104] <= 3'b000;
      memory_array[8105] <= 3'b101;
      memory_array[8106] <= 3'b000;
      memory_array[8107] <= 3'b101;
      memory_array[8108] <= 3'b000;
      memory_array[8109] <= 3'b000;
      memory_array[8110] <= 3'b101;
      memory_array[8111] <= 3'b101;
      memory_array[8112] <= 3'b101;
      memory_array[8113] <= 3'b101;
      memory_array[8114] <= 3'b000;
      memory_array[8115] <= 3'b101;
      memory_array[8116] <= 3'b000;
      memory_array[8117] <= 3'b000;
      memory_array[8118] <= 3'b101;
      memory_array[8119] <= 3'b101;
      memory_array[8120] <= 3'b000;
      memory_array[8121] <= 3'b101;
      memory_array[8122] <= 3'b101;
      memory_array[8123] <= 3'b000;
      memory_array[8124] <= 3'b101;
      memory_array[8125] <= 3'b101;
      memory_array[8126] <= 3'b101;
      memory_array[8127] <= 3'b101;
      memory_array[8128] <= 3'b000;
      memory_array[8129] <= 3'b101;
      memory_array[8130] <= 3'b101;
      memory_array[8131] <= 3'b101;
      memory_array[8132] <= 3'b000;
      memory_array[8133] <= 3'b101;
      memory_array[8134] <= 3'b101;
      memory_array[8135] <= 3'b101;
      memory_array[8136] <= 3'b101;
      memory_array[8137] <= 3'b000;
      memory_array[8138] <= 3'b101;
      memory_array[8139] <= 3'b000;
      memory_array[8140] <= 3'b101;
      memory_array[8141] <= 3'b101;
      memory_array[8142] <= 3'b101;
      memory_array[8143] <= 3'b000;
      memory_array[8144] <= 3'b101;
      memory_array[8145] <= 3'b101;
      memory_array[8146] <= 3'b101;
      memory_array[8147] <= 3'b101;
      memory_array[8148] <= 3'b101;
      memory_array[8149] <= 3'b000;
      memory_array[8150] <= 3'b101;
      memory_array[8151] <= 3'b101;
      memory_array[8152] <= 3'b101;
      memory_array[8153] <= 3'b000;
      memory_array[8154] <= 3'b101;
      memory_array[8155] <= 3'b101;
      memory_array[8156] <= 3'b000;
      memory_array[8157] <= 3'b111;
      memory_array[8158] <= 3'b111;
      memory_array[8159] <= 3'b111;
      memory_array[8160] <= 3'b111;
      memory_array[8161] <= 3'b111;
      memory_array[8162] <= 3'b000;
      memory_array[8163] <= 3'b000;
      memory_array[8164] <= 3'b000;
      memory_array[8165] <= 3'b110;
      memory_array[8166] <= 3'b110;
      memory_array[8167] <= 3'b110;
      memory_array[8168] <= 3'b000;
      memory_array[8169] <= 3'b000;
      memory_array[8170] <= 3'b000;
      memory_array[8171] <= 3'b000;
      memory_array[8172] <= 3'b000;
      memory_array[8173] <= 3'b101;
      memory_array[8174] <= 3'b000;
      memory_array[8175] <= 3'b000;
      memory_array[8176] <= 3'b110;
      memory_array[8177] <= 3'b110;
      memory_array[8178] <= 3'b000;
      memory_array[8179] <= 3'b000;
      memory_array[8180] <= 3'b110;
      memory_array[8181] <= 3'b110;
      memory_array[8182] <= 3'b110;
      memory_array[8183] <= 3'b000;
      memory_array[8184] <= 3'b000;
      memory_array[8185] <= 3'b110;
      memory_array[8186] <= 3'b101;
      memory_array[8187] <= 3'b110;
      memory_array[8188] <= 3'b000;
      memory_array[8189] <= 3'b000;
      memory_array[8190] <= 3'b000;
      memory_array[8191] <= 3'b101;
      memory_array[8192] <= 3'b101;
      memory_array[8193] <= 3'b101;
      memory_array[8194] <= 3'b101;
      memory_array[8195] <= 3'b101;
      memory_array[8196] <= 3'b101;
      memory_array[8197] <= 3'b101;
      memory_array[8198] <= 3'b101;
      memory_array[8199] <= 3'b101;
      memory_array[8200] <= 3'b101;
      memory_array[8201] <= 3'b101;
      memory_array[8202] <= 3'b101;
      memory_array[8203] <= 3'b101;
      memory_array[8204] <= 3'b101;
      memory_array[8205] <= 3'b101;
      memory_array[8206] <= 3'b101;
      memory_array[8207] <= 3'b101;
      memory_array[8208] <= 3'b101;
      memory_array[8209] <= 3'b000;
      memory_array[8210] <= 3'b000;
      memory_array[8211] <= 3'b110;
      memory_array[8212] <= 3'b000;
      memory_array[8213] <= 3'b000;
      memory_array[8214] <= 3'b000;
      memory_array[8215] <= 3'b110;
      memory_array[8216] <= 3'b110;
      memory_array[8217] <= 3'b110;
      memory_array[8218] <= 3'b000;
      memory_array[8219] <= 3'b000;
      memory_array[8220] <= 3'b110;
      memory_array[8221] <= 3'b110;
      memory_array[8222] <= 3'b110;
      memory_array[8223] <= 3'b000;
      memory_array[8224] <= 3'b000;
      memory_array[8225] <= 3'b110;
      memory_array[8226] <= 3'b000;
      memory_array[8227] <= 3'b000;
      memory_array[8228] <= 3'b000;
      memory_array[8229] <= 3'b000;
      memory_array[8230] <= 3'b110;
      memory_array[8231] <= 3'b110;
      memory_array[8232] <= 3'b110;
      memory_array[8233] <= 3'b000;
      memory_array[8234] <= 3'b000;
      memory_array[8235] <= 3'b110;
      memory_array[8236] <= 3'b000;
      memory_array[8237] <= 3'b111;
      memory_array[8238] <= 3'b111;
      memory_array[8239] <= 3'b111;
      memory_array[8240] <= 3'b111;
      memory_array[8241] <= 3'b101;
      memory_array[8242] <= 3'b101;
      memory_array[8243] <= 3'b101;
      memory_array[8244] <= 3'b101;
      memory_array[8245] <= 3'b101;
      memory_array[8246] <= 3'b101;
      memory_array[8247] <= 3'b101;
      memory_array[8248] <= 3'b000;
      memory_array[8249] <= 3'b000;
      memory_array[8250] <= 3'b101;
      memory_array[8251] <= 3'b101;
      memory_array[8252] <= 3'b101;
      memory_array[8253] <= 3'b000;
      memory_array[8254] <= 3'b101;
      memory_array[8255] <= 3'b101;
      memory_array[8256] <= 3'b111;
      memory_array[8257] <= 3'b101;
      memory_array[8258] <= 3'b101;
      memory_array[8259] <= 3'b101;
      memory_array[8260] <= 3'b101;
      memory_array[8261] <= 3'b101;
      memory_array[8262] <= 3'b000;
      memory_array[8263] <= 3'b101;
      memory_array[8264] <= 3'b101;
      memory_array[8265] <= 3'b101;
      memory_array[8266] <= 3'b101;
      memory_array[8267] <= 3'b000;
      memory_array[8268] <= 3'b101;
      memory_array[8269] <= 3'b101;
      memory_array[8270] <= 3'b101;
      memory_array[8271] <= 3'b101;
      memory_array[8272] <= 3'b101;
      memory_array[8273] <= 3'b101;
      memory_array[8274] <= 3'b111;
      memory_array[8275] <= 3'b101;
      memory_array[8276] <= 3'b000;
      memory_array[8277] <= 3'b101;
      memory_array[8278] <= 3'b101;
      memory_array[8279] <= 3'b101;
      memory_array[8280] <= 3'b101;
      memory_array[8281] <= 3'b111;
      memory_array[8282] <= 3'b111;
      memory_array[8283] <= 3'b111;
      memory_array[8284] <= 3'b111;
      memory_array[8285] <= 3'b111;
      memory_array[8286] <= 3'b111;
      memory_array[8287] <= 3'b111;
      memory_array[8288] <= 3'b111;
      memory_array[8289] <= 3'b000;
      memory_array[8290] <= 3'b101;
      memory_array[8291] <= 3'b111;
      memory_array[8292] <= 3'b101;
      memory_array[8293] <= 3'b111;
      memory_array[8294] <= 3'b000;
      memory_array[8295] <= 3'b101;
      memory_array[8296] <= 3'b000;
      memory_array[8297] <= 3'b111;
      memory_array[8298] <= 3'b111;
      memory_array[8299] <= 3'b000;
      memory_array[8300] <= 3'b101;
      memory_array[8301] <= 3'b111;
      memory_array[8302] <= 3'b111;
      memory_array[8303] <= 3'b000;
      memory_array[8304] <= 3'b101;
      memory_array[8305] <= 3'b101;
      memory_array[8306] <= 3'b000;
      memory_array[8307] <= 3'b101;
      memory_array[8308] <= 3'b101;
      memory_array[8309] <= 3'b101;
      memory_array[8310] <= 3'b101;
      memory_array[8311] <= 3'b101;
      memory_array[8312] <= 3'b000;
      memory_array[8313] <= 3'b000;
      memory_array[8314] <= 3'b101;
      memory_array[8315] <= 3'b101;
      memory_array[8316] <= 3'b101;
      memory_array[8317] <= 3'b101;
      memory_array[8318] <= 3'b101;
      memory_array[8319] <= 3'b101;
      memory_array[8320] <= 3'b101;
      memory_array[8321] <= 3'b101;
      memory_array[8322] <= 3'b101;
      memory_array[8323] <= 3'b101;
      memory_array[8324] <= 3'b101;
      memory_array[8325] <= 3'b101;
      memory_array[8326] <= 3'b000;
      memory_array[8327] <= 3'b101;
      memory_array[8328] <= 3'b101;
      memory_array[8329] <= 3'b101;
      memory_array[8330] <= 3'b101;
      memory_array[8331] <= 3'b111;
      memory_array[8332] <= 3'b101;
      memory_array[8333] <= 3'b101;
      memory_array[8334] <= 3'b101;
      memory_array[8335] <= 3'b101;
      memory_array[8336] <= 3'b101;
      memory_array[8337] <= 3'b101;
      memory_array[8338] <= 3'b101;
      memory_array[8339] <= 3'b101;
      memory_array[8340] <= 3'b101;
      memory_array[8341] <= 3'b101;
      memory_array[8342] <= 3'b101;
      memory_array[8343] <= 3'b101;
      memory_array[8344] <= 3'b101;
      memory_array[8345] <= 3'b101;
      memory_array[8346] <= 3'b000;
      memory_array[8347] <= 3'b101;
      memory_array[8348] <= 3'b101;
      memory_array[8349] <= 3'b101;
      memory_array[8350] <= 3'b000;
      memory_array[8351] <= 3'b000;
      memory_array[8352] <= 3'b000;
      memory_array[8353] <= 3'b101;
      memory_array[8354] <= 3'b101;
      memory_array[8355] <= 3'b101;
      memory_array[8356] <= 3'b101;
      memory_array[8357] <= 3'b000;
      memory_array[8358] <= 3'b101;
      memory_array[8359] <= 3'b111;
      memory_array[8360] <= 3'b111;
      memory_array[8361] <= 3'b111;
      memory_array[8362] <= 3'b101;
      memory_array[8363] <= 3'b000;
      memory_array[8364] <= 3'b000;
      memory_array[8365] <= 3'b110;
      memory_array[8366] <= 3'b110;
      memory_array[8367] <= 3'b110;
      memory_array[8368] <= 3'b000;
      memory_array[8369] <= 3'b000;
      memory_array[8370] <= 3'b110;
      memory_array[8371] <= 3'b110;
      memory_array[8372] <= 3'b000;
      memory_array[8373] <= 3'b000;
      memory_array[8374] <= 3'b000;
      memory_array[8375] <= 3'b110;
      memory_array[8376] <= 3'b110;
      memory_array[8377] <= 3'b110;
      memory_array[8378] <= 3'b000;
      memory_array[8379] <= 3'b000;
      memory_array[8380] <= 3'b110;
      memory_array[8381] <= 3'b110;
      memory_array[8382] <= 3'b110;
      memory_array[8383] <= 3'b000;
      memory_array[8384] <= 3'b000;
      memory_array[8385] <= 3'b110;
      memory_array[8386] <= 3'b110;
      memory_array[8387] <= 3'b110;
      memory_array[8388] <= 3'b000;
      memory_array[8389] <= 3'b000;
      memory_array[8390] <= 3'b000;
      memory_array[8391] <= 3'b101;
      memory_array[8392] <= 3'b101;
      memory_array[8393] <= 3'b101;
      memory_array[8394] <= 3'b101;
      memory_array[8395] <= 3'b101;
      memory_array[8396] <= 3'b101;
      memory_array[8397] <= 3'b101;
      memory_array[8398] <= 3'b101;
      memory_array[8399] <= 3'b101;
      memory_array[8400] <= 3'b101;
      memory_array[8401] <= 3'b101;
      memory_array[8402] <= 3'b101;
      memory_array[8403] <= 3'b111;
      memory_array[8404] <= 3'b111;
      memory_array[8405] <= 3'b101;
      memory_array[8406] <= 3'b101;
      memory_array[8407] <= 3'b101;
      memory_array[8408] <= 3'b101;
      memory_array[8409] <= 3'b000;
      memory_array[8410] <= 3'b000;
      memory_array[8411] <= 3'b000;
      memory_array[8412] <= 3'b000;
      memory_array[8413] <= 3'b110;
      memory_array[8414] <= 3'b110;
      memory_array[8415] <= 3'b000;
      memory_array[8416] <= 3'b000;
      memory_array[8417] <= 3'b000;
      memory_array[8418] <= 3'b101;
      memory_array[8419] <= 3'b000;
      memory_array[8420] <= 3'b000;
      memory_array[8421] <= 3'b101;
      memory_array[8422] <= 3'b000;
      memory_array[8423] <= 3'b110;
      memory_array[8424] <= 3'b110;
      memory_array[8425] <= 3'b000;
      memory_array[8426] <= 3'b000;
      memory_array[8427] <= 3'b000;
      memory_array[8428] <= 3'b110;
      memory_array[8429] <= 3'b110;
      memory_array[8430] <= 3'b000;
      memory_array[8431] <= 3'b000;
      memory_array[8432] <= 3'b000;
      memory_array[8433] <= 3'b110;
      memory_array[8434] <= 3'b110;
      memory_array[8435] <= 3'b000;
      memory_array[8436] <= 3'b101;
      memory_array[8437] <= 3'b111;
      memory_array[8438] <= 3'b111;
      memory_array[8439] <= 3'b111;
      memory_array[8440] <= 3'b111;
      memory_array[8441] <= 3'b000;
      memory_array[8442] <= 3'b101;
      memory_array[8443] <= 3'b101;
      memory_array[8444] <= 3'b101;
      memory_array[8445] <= 3'b000;
      memory_array[8446] <= 3'b101;
      memory_array[8447] <= 3'b101;
      memory_array[8448] <= 3'b101;
      memory_array[8449] <= 3'b101;
      memory_array[8450] <= 3'b000;
      memory_array[8451] <= 3'b101;
      memory_array[8452] <= 3'b101;
      memory_array[8453] <= 3'b000;
      memory_array[8454] <= 3'b101;
      memory_array[8455] <= 3'b101;
      memory_array[8456] <= 3'b111;
      memory_array[8457] <= 3'b000;
      memory_array[8458] <= 3'b000;
      memory_array[8459] <= 3'b000;
      memory_array[8460] <= 3'b101;
      memory_array[8461] <= 3'b101;
      memory_array[8462] <= 3'b101;
      memory_array[8463] <= 3'b101;
      memory_array[8464] <= 3'b101;
      memory_array[8465] <= 3'b101;
      memory_array[8466] <= 3'b101;
      memory_array[8467] <= 3'b101;
      memory_array[8468] <= 3'b101;
      memory_array[8469] <= 3'b101;
      memory_array[8470] <= 3'b000;
      memory_array[8471] <= 3'b101;
      memory_array[8472] <= 3'b101;
      memory_array[8473] <= 3'b101;
      memory_array[8474] <= 3'b111;
      memory_array[8475] <= 3'b111;
      memory_array[8476] <= 3'b000;
      memory_array[8477] <= 3'b000;
      memory_array[8478] <= 3'b101;
      memory_array[8479] <= 3'b000;
      memory_array[8480] <= 3'b101;
      memory_array[8481] <= 3'b111;
      memory_array[8482] <= 3'b111;
      memory_array[8483] <= 3'b111;
      memory_array[8484] <= 3'b111;
      memory_array[8485] <= 3'b111;
      memory_array[8486] <= 3'b111;
      memory_array[8487] <= 3'b111;
      memory_array[8488] <= 3'b111;
      memory_array[8489] <= 3'b000;
      memory_array[8490] <= 3'b000;
      memory_array[8491] <= 3'b111;
      memory_array[8492] <= 3'b000;
      memory_array[8493] <= 3'b111;
      memory_array[8494] <= 3'b000;
      memory_array[8495] <= 3'b101;
      memory_array[8496] <= 3'b000;
      memory_array[8497] <= 3'b000;
      memory_array[8498] <= 3'b101;
      memory_array[8499] <= 3'b101;
      memory_array[8500] <= 3'b101;
      memory_array[8501] <= 3'b111;
      memory_array[8502] <= 3'b111;
      memory_array[8503] <= 3'b000;
      memory_array[8504] <= 3'b101;
      memory_array[8505] <= 3'b101;
      memory_array[8506] <= 3'b101;
      memory_array[8507] <= 3'b101;
      memory_array[8508] <= 3'b101;
      memory_array[8509] <= 3'b101;
      memory_array[8510] <= 3'b101;
      memory_array[8511] <= 3'b000;
      memory_array[8512] <= 3'b101;
      memory_array[8513] <= 3'b101;
      memory_array[8514] <= 3'b000;
      memory_array[8515] <= 3'b101;
      memory_array[8516] <= 3'b101;
      memory_array[8517] <= 3'b101;
      memory_array[8518] <= 3'b101;
      memory_array[8519] <= 3'b101;
      memory_array[8520] <= 3'b000;
      memory_array[8521] <= 3'b101;
      memory_array[8522] <= 3'b101;
      memory_array[8523] <= 3'b101;
      memory_array[8524] <= 3'b101;
      memory_array[8525] <= 3'b101;
      memory_array[8526] <= 3'b101;
      memory_array[8527] <= 3'b101;
      memory_array[8528] <= 3'b101;
      memory_array[8529] <= 3'b000;
      memory_array[8530] <= 3'b101;
      memory_array[8531] <= 3'b111;
      memory_array[8532] <= 3'b000;
      memory_array[8533] <= 3'b101;
      memory_array[8534] <= 3'b101;
      memory_array[8535] <= 3'b101;
      memory_array[8536] <= 3'b101;
      memory_array[8537] <= 3'b101;
      memory_array[8538] <= 3'b101;
      memory_array[8539] <= 3'b101;
      memory_array[8540] <= 3'b000;
      memory_array[8541] <= 3'b000;
      memory_array[8542] <= 3'b101;
      memory_array[8543] <= 3'b101;
      memory_array[8544] <= 3'b101;
      memory_array[8545] <= 3'b101;
      memory_array[8546] <= 3'b000;
      memory_array[8547] <= 3'b000;
      memory_array[8548] <= 3'b101;
      memory_array[8549] <= 3'b000;
      memory_array[8550] <= 3'b101;
      memory_array[8551] <= 3'b101;
      memory_array[8552] <= 3'b000;
      memory_array[8553] <= 3'b101;
      memory_array[8554] <= 3'b000;
      memory_array[8555] <= 3'b101;
      memory_array[8556] <= 3'b101;
      memory_array[8557] <= 3'b000;
      memory_array[8558] <= 3'b000;
      memory_array[8559] <= 3'b111;
      memory_array[8560] <= 3'b111;
      memory_array[8561] <= 3'b111;
      memory_array[8562] <= 3'b111;
      memory_array[8563] <= 3'b101;
      memory_array[8564] <= 3'b110;
      memory_array[8565] <= 3'b000;
      memory_array[8566] <= 3'b000;
      memory_array[8567] <= 3'b000;
      memory_array[8568] <= 3'b110;
      memory_array[8569] <= 3'b110;
      memory_array[8570] <= 3'b000;
      memory_array[8571] <= 3'b000;
      memory_array[8572] <= 3'b000;
      memory_array[8573] <= 3'b110;
      memory_array[8574] <= 3'b110;
      memory_array[8575] <= 3'b000;
      memory_array[8576] <= 3'b000;
      memory_array[8577] <= 3'b000;
      memory_array[8578] <= 3'b101;
      memory_array[8579] <= 3'b110;
      memory_array[8580] <= 3'b000;
      memory_array[8581] <= 3'b101;
      memory_array[8582] <= 3'b000;
      memory_array[8583] <= 3'b110;
      memory_array[8584] <= 3'b110;
      memory_array[8585] <= 3'b000;
      memory_array[8586] <= 3'b000;
      memory_array[8587] <= 3'b000;
      memory_array[8588] <= 3'b110;
      memory_array[8589] <= 3'b000;
      memory_array[8590] <= 3'b000;
      memory_array[8591] <= 3'b101;
      memory_array[8592] <= 3'b101;
      memory_array[8593] <= 3'b101;
      memory_array[8594] <= 3'b101;
      memory_array[8595] <= 3'b111;
      memory_array[8596] <= 3'b111;
      memory_array[8597] <= 3'b101;
      memory_array[8598] <= 3'b101;
      memory_array[8599] <= 3'b101;
      memory_array[8600] <= 3'b101;
      memory_array[8601] <= 3'b101;
      memory_array[8602] <= 3'b110;
      memory_array[8603] <= 3'b101;
      memory_array[8604] <= 3'b101;
      memory_array[8605] <= 3'b110;
      memory_array[8606] <= 3'b101;
      memory_array[8607] <= 3'b101;
      memory_array[8608] <= 3'b101;
      memory_array[8609] <= 3'b000;
      memory_array[8610] <= 3'b000;
      memory_array[8611] <= 3'b110;
      memory_array[8612] <= 3'b110;
      memory_array[8613] <= 3'b000;
      memory_array[8614] <= 3'b000;
      memory_array[8615] <= 3'b110;
      memory_array[8616] <= 3'b110;
      memory_array[8617] <= 3'b000;
      memory_array[8618] <= 3'b000;
      memory_array[8619] <= 3'b101;
      memory_array[8620] <= 3'b101;
      memory_array[8621] <= 3'b000;
      memory_array[8622] <= 3'b110;
      memory_array[8623] <= 3'b000;
      memory_array[8624] <= 3'b000;
      memory_array[8625] <= 3'b110;
      memory_array[8626] <= 3'b000;
      memory_array[8627] <= 3'b110;
      memory_array[8628] <= 3'b000;
      memory_array[8629] <= 3'b000;
      memory_array[8630] <= 3'b101;
      memory_array[8631] <= 3'b000;
      memory_array[8632] <= 3'b110;
      memory_array[8633] <= 3'b000;
      memory_array[8634] <= 3'b000;
      memory_array[8635] <= 3'b000;
      memory_array[8636] <= 3'b111;
      memory_array[8637] <= 3'b111;
      memory_array[8638] <= 3'b111;
      memory_array[8639] <= 3'b111;
      memory_array[8640] <= 3'b111;
      memory_array[8641] <= 3'b000;
      memory_array[8642] <= 3'b101;
      memory_array[8643] <= 3'b101;
      memory_array[8644] <= 3'b101;
      memory_array[8645] <= 3'b101;
      memory_array[8646] <= 3'b101;
      memory_array[8647] <= 3'b101;
      memory_array[8648] <= 3'b101;
      memory_array[8649] <= 3'b101;
      memory_array[8650] <= 3'b101;
      memory_array[8651] <= 3'b000;
      memory_array[8652] <= 3'b101;
      memory_array[8653] <= 3'b101;
      memory_array[8654] <= 3'b101;
      memory_array[8655] <= 3'b000;
      memory_array[8656] <= 3'b101;
      memory_array[8657] <= 3'b000;
      memory_array[8658] <= 3'b000;
      memory_array[8659] <= 3'b101;
      memory_array[8660] <= 3'b101;
      memory_array[8661] <= 3'b101;
      memory_array[8662] <= 3'b101;
      memory_array[8663] <= 3'b101;
      memory_array[8664] <= 3'b101;
      memory_array[8665] <= 3'b101;
      memory_array[8666] <= 3'b101;
      memory_array[8667] <= 3'b000;
      memory_array[8668] <= 3'b101;
      memory_array[8669] <= 3'b101;
      memory_array[8670] <= 3'b101;
      memory_array[8671] <= 3'b101;
      memory_array[8672] <= 3'b101;
      memory_array[8673] <= 3'b000;
      memory_array[8674] <= 3'b111;
      memory_array[8675] <= 3'b111;
      memory_array[8676] <= 3'b101;
      memory_array[8677] <= 3'b101;
      memory_array[8678] <= 3'b000;
      memory_array[8679] <= 3'b101;
      memory_array[8680] <= 3'b111;
      memory_array[8681] <= 3'b111;
      memory_array[8682] <= 3'b111;
      memory_array[8683] <= 3'b111;
      memory_array[8684] <= 3'b111;
      memory_array[8685] <= 3'b111;
      memory_array[8686] <= 3'b111;
      memory_array[8687] <= 3'b111;
      memory_array[8688] <= 3'b111;
      memory_array[8689] <= 3'b101;
      memory_array[8690] <= 3'b000;
      memory_array[8691] <= 3'b101;
      memory_array[8692] <= 3'b101;
      memory_array[8693] <= 3'b111;
      memory_array[8694] <= 3'b000;
      memory_array[8695] <= 3'b101;
      memory_array[8696] <= 3'b000;
      memory_array[8697] <= 3'b111;
      memory_array[8698] <= 3'b000;
      memory_array[8699] <= 3'b101;
      memory_array[8700] <= 3'b111;
      memory_array[8701] <= 3'b111;
      memory_array[8702] <= 3'b111;
      memory_array[8703] <= 3'b000;
      memory_array[8704] <= 3'b000;
      memory_array[8705] <= 3'b101;
      memory_array[8706] <= 3'b101;
      memory_array[8707] <= 3'b000;
      memory_array[8708] <= 3'b101;
      memory_array[8709] <= 3'b101;
      memory_array[8710] <= 3'b101;
      memory_array[8711] <= 3'b101;
      memory_array[8712] <= 3'b101;
      memory_array[8713] <= 3'b101;
      memory_array[8714] <= 3'b101;
      memory_array[8715] <= 3'b101;
      memory_array[8716] <= 3'b101;
      memory_array[8717] <= 3'b101;
      memory_array[8718] <= 3'b101;
      memory_array[8719] <= 3'b101;
      memory_array[8720] <= 3'b101;
      memory_array[8721] <= 3'b000;
      memory_array[8722] <= 3'b101;
      memory_array[8723] <= 3'b101;
      memory_array[8724] <= 3'b101;
      memory_array[8725] <= 3'b101;
      memory_array[8726] <= 3'b000;
      memory_array[8727] <= 3'b101;
      memory_array[8728] <= 3'b101;
      memory_array[8729] <= 3'b101;
      memory_array[8730] <= 3'b101;
      memory_array[8731] <= 3'b101;
      memory_array[8732] <= 3'b101;
      memory_array[8733] <= 3'b101;
      memory_array[8734] <= 3'b101;
      memory_array[8735] <= 3'b101;
      memory_array[8736] <= 3'b101;
      memory_array[8737] <= 3'b101;
      memory_array[8738] <= 3'b101;
      memory_array[8739] <= 3'b101;
      memory_array[8740] <= 3'b101;
      memory_array[8741] <= 3'b000;
      memory_array[8742] <= 3'b101;
      memory_array[8743] <= 3'b101;
      memory_array[8744] <= 3'b000;
      memory_array[8745] <= 3'b101;
      memory_array[8746] <= 3'b101;
      memory_array[8747] <= 3'b000;
      memory_array[8748] <= 3'b000;
      memory_array[8749] <= 3'b101;
      memory_array[8750] <= 3'b101;
      memory_array[8751] <= 3'b101;
      memory_array[8752] <= 3'b101;
      memory_array[8753] <= 3'b101;
      memory_array[8754] <= 3'b101;
      memory_array[8755] <= 3'b101;
      memory_array[8756] <= 3'b101;
      memory_array[8757] <= 3'b101;
      memory_array[8758] <= 3'b000;
      memory_array[8759] <= 3'b111;
      memory_array[8760] <= 3'b111;
      memory_array[8761] <= 3'b111;
      memory_array[8762] <= 3'b111;
      memory_array[8763] <= 3'b111;
      memory_array[8764] <= 3'b000;
      memory_array[8765] <= 3'b110;
      memory_array[8766] <= 3'b110;
      memory_array[8767] <= 3'b110;
      memory_array[8768] <= 3'b000;
      memory_array[8769] <= 3'b101;
      memory_array[8770] <= 3'b000;
      memory_array[8771] <= 3'b110;
      memory_array[8772] <= 3'b000;
      memory_array[8773] <= 3'b000;
      memory_array[8774] <= 3'b000;
      memory_array[8775] <= 3'b110;
      memory_array[8776] <= 3'b110;
      memory_array[8777] <= 3'b110;
      memory_array[8778] <= 3'b000;
      memory_array[8779] <= 3'b101;
      memory_array[8780] <= 3'b101;
      memory_array[8781] <= 3'b000;
      memory_array[8782] <= 3'b110;
      memory_array[8783] <= 3'b000;
      memory_array[8784] <= 3'b000;
      memory_array[8785] <= 3'b110;
      memory_array[8786] <= 3'b110;
      memory_array[8787] <= 3'b110;
      memory_array[8788] <= 3'b000;
      memory_array[8789] <= 3'b000;
      memory_array[8790] <= 3'b000;
      memory_array[8791] <= 3'b101;
      memory_array[8792] <= 3'b101;
      memory_array[8793] <= 3'b101;
      memory_array[8794] <= 3'b000;
      memory_array[8795] <= 3'b101;
      memory_array[8796] <= 3'b101;
      memory_array[8797] <= 3'b110;
      memory_array[8798] <= 3'b101;
      memory_array[8799] <= 3'b101;
      memory_array[8800] <= 3'b110;
      memory_array[8801] <= 3'b110;
      memory_array[8802] <= 3'b110;
      memory_array[8803] <= 3'b000;
      memory_array[8804] <= 3'b000;
      memory_array[8805] <= 3'b110;
      memory_array[8806] <= 3'b110;
      memory_array[8807] <= 3'b101;
      memory_array[8808] <= 3'b101;
      memory_array[8809] <= 3'b000;
      memory_array[8810] <= 3'b000;
      memory_array[8811] <= 3'b110;
      memory_array[8812] <= 3'b110;
      memory_array[8813] <= 3'b000;
      memory_array[8814] <= 3'b000;
      memory_array[8815] <= 3'b110;
      memory_array[8816] <= 3'b110;
      memory_array[8817] <= 3'b110;
      memory_array[8818] <= 3'b000;
      memory_array[8819] <= 3'b000;
      memory_array[8820] <= 3'b000;
      memory_array[8821] <= 3'b000;
      memory_array[8822] <= 3'b000;
      memory_array[8823] <= 3'b101;
      memory_array[8824] <= 3'b101;
      memory_array[8825] <= 3'b101;
      memory_array[8826] <= 3'b110;
      memory_array[8827] <= 3'b110;
      memory_array[8828] <= 3'b000;
      memory_array[8829] <= 3'b000;
      memory_array[8830] <= 3'b000;
      memory_array[8831] <= 3'b110;
      memory_array[8832] <= 3'b110;
      memory_array[8833] <= 3'b000;
      memory_array[8834] <= 3'b000;
      memory_array[8835] <= 3'b000;
      memory_array[8836] <= 3'b111;
      memory_array[8837] <= 3'b111;
      memory_array[8838] <= 3'b111;
      memory_array[8839] <= 3'b111;
      memory_array[8840] <= 3'b101;
      memory_array[8841] <= 3'b101;
      memory_array[8842] <= 3'b101;
      memory_array[8843] <= 3'b101;
      memory_array[8844] <= 3'b101;
      memory_array[8845] <= 3'b101;
      memory_array[8846] <= 3'b101;
      memory_array[8847] <= 3'b101;
      memory_array[8848] <= 3'b101;
      memory_array[8849] <= 3'b101;
      memory_array[8850] <= 3'b101;
      memory_array[8851] <= 3'b101;
      memory_array[8852] <= 3'b101;
      memory_array[8853] <= 3'b101;
      memory_array[8854] <= 3'b000;
      memory_array[8855] <= 3'b101;
      memory_array[8856] <= 3'b101;
      memory_array[8857] <= 3'b101;
      memory_array[8858] <= 3'b101;
      memory_array[8859] <= 3'b101;
      memory_array[8860] <= 3'b000;
      memory_array[8861] <= 3'b101;
      memory_array[8862] <= 3'b101;
      memory_array[8863] <= 3'b101;
      memory_array[8864] <= 3'b101;
      memory_array[8865] <= 3'b101;
      memory_array[8866] <= 3'b101;
      memory_array[8867] <= 3'b101;
      memory_array[8868] <= 3'b000;
      memory_array[8869] <= 3'b101;
      memory_array[8870] <= 3'b000;
      memory_array[8871] <= 3'b101;
      memory_array[8872] <= 3'b101;
      memory_array[8873] <= 3'b101;
      memory_array[8874] <= 3'b110;
      memory_array[8875] <= 3'b101;
      memory_array[8876] <= 3'b101;
      memory_array[8877] <= 3'b101;
      memory_array[8878] <= 3'b000;
      memory_array[8879] <= 3'b111;
      memory_array[8880] <= 3'b111;
      memory_array[8881] <= 3'b111;
      memory_array[8882] <= 3'b111;
      memory_array[8883] <= 3'b111;
      memory_array[8884] <= 3'b111;
      memory_array[8885] <= 3'b111;
      memory_array[8886] <= 3'b111;
      memory_array[8887] <= 3'b111;
      memory_array[8888] <= 3'b111;
      memory_array[8889] <= 3'b101;
      memory_array[8890] <= 3'b101;
      memory_array[8891] <= 3'b000;
      memory_array[8892] <= 3'b101;
      memory_array[8893] <= 3'b111;
      memory_array[8894] <= 3'b000;
      memory_array[8895] <= 3'b101;
      memory_array[8896] <= 3'b101;
      memory_array[8897] <= 3'b101;
      memory_array[8898] <= 3'b111;
      memory_array[8899] <= 3'b111;
      memory_array[8900] <= 3'b101;
      memory_array[8901] <= 3'b111;
      memory_array[8902] <= 3'b111;
      memory_array[8903] <= 3'b000;
      memory_array[8904] <= 3'b101;
      memory_array[8905] <= 3'b101;
      memory_array[8906] <= 3'b000;
      memory_array[8907] <= 3'b101;
      memory_array[8908] <= 3'b101;
      memory_array[8909] <= 3'b101;
      memory_array[8910] <= 3'b101;
      memory_array[8911] <= 3'b101;
      memory_array[8912] <= 3'b101;
      memory_array[8913] <= 3'b101;
      memory_array[8914] <= 3'b101;
      memory_array[8915] <= 3'b101;
      memory_array[8916] <= 3'b101;
      memory_array[8917] <= 3'b101;
      memory_array[8918] <= 3'b101;
      memory_array[8919] <= 3'b101;
      memory_array[8920] <= 3'b101;
      memory_array[8921] <= 3'b000;
      memory_array[8922] <= 3'b101;
      memory_array[8923] <= 3'b101;
      memory_array[8924] <= 3'b101;
      memory_array[8925] <= 3'b000;
      memory_array[8926] <= 3'b101;
      memory_array[8927] <= 3'b101;
      memory_array[8928] <= 3'b101;
      memory_array[8929] <= 3'b000;
      memory_array[8930] <= 3'b101;
      memory_array[8931] <= 3'b000;
      memory_array[8932] <= 3'b101;
      memory_array[8933] <= 3'b101;
      memory_array[8934] <= 3'b101;
      memory_array[8935] <= 3'b101;
      memory_array[8936] <= 3'b101;
      memory_array[8937] <= 3'b101;
      memory_array[8938] <= 3'b101;
      memory_array[8939] <= 3'b000;
      memory_array[8940] <= 3'b101;
      memory_array[8941] <= 3'b101;
      memory_array[8942] <= 3'b101;
      memory_array[8943] <= 3'b101;
      memory_array[8944] <= 3'b101;
      memory_array[8945] <= 3'b000;
      memory_array[8946] <= 3'b101;
      memory_array[8947] <= 3'b101;
      memory_array[8948] <= 3'b101;
      memory_array[8949] <= 3'b101;
      memory_array[8950] <= 3'b101;
      memory_array[8951] <= 3'b101;
      memory_array[8952] <= 3'b101;
      memory_array[8953] <= 3'b101;
      memory_array[8954] <= 3'b101;
      memory_array[8955] <= 3'b101;
      memory_array[8956] <= 3'b101;
      memory_array[8957] <= 3'b000;
      memory_array[8958] <= 3'b101;
      memory_array[8959] <= 3'b101;
      memory_array[8960] <= 3'b111;
      memory_array[8961] <= 3'b111;
      memory_array[8962] <= 3'b111;
      memory_array[8963] <= 3'b111;
      memory_array[8964] <= 3'b000;
      memory_array[8965] <= 3'b000;
      memory_array[8966] <= 3'b110;
      memory_array[8967] <= 3'b110;
      memory_array[8968] <= 3'b000;
      memory_array[8969] <= 3'b000;
      memory_array[8970] <= 3'b000;
      memory_array[8971] <= 3'b110;
      memory_array[8972] <= 3'b110;
      memory_array[8973] <= 3'b000;
      memory_array[8974] <= 3'b101;
      memory_array[8975] <= 3'b101;
      memory_array[8976] <= 3'b101;
      memory_array[8977] <= 3'b000;
      memory_array[8978] <= 3'b000;
      memory_array[8979] <= 3'b000;
      memory_array[8980] <= 3'b110;
      memory_array[8981] <= 3'b110;
      memory_array[8982] <= 3'b110;
      memory_array[8983] <= 3'b000;
      memory_array[8984] <= 3'b000;
      memory_array[8985] <= 3'b110;
      memory_array[8986] <= 3'b110;
      memory_array[8987] <= 3'b110;
      memory_array[8988] <= 3'b000;
      memory_array[8989] <= 3'b000;
      memory_array[8990] <= 3'b000;
      memory_array[8991] <= 3'b101;
      memory_array[8992] <= 3'b110;
      memory_array[8993] <= 3'b000;
      memory_array[8994] <= 3'b000;
      memory_array[8995] <= 3'b110;
      memory_array[8996] <= 3'b110;
      memory_array[8997] <= 3'b110;
      memory_array[8998] <= 3'b000;
      memory_array[8999] <= 3'b101;
      memory_array[9000] <= 3'b000;
      memory_array[9001] <= 3'b000;
      memory_array[9002] <= 3'b000;
      memory_array[9003] <= 3'b110;
      memory_array[9004] <= 3'b110;
      memory_array[9005] <= 3'b000;
      memory_array[9006] <= 3'b000;
      memory_array[9007] <= 3'b000;
      memory_array[9008] <= 3'b101;
      memory_array[9009] <= 3'b000;
      memory_array[9010] <= 3'b000;
      memory_array[9011] <= 3'b000;
      memory_array[9012] <= 3'b000;
      memory_array[9013] <= 3'b110;
      memory_array[9014] <= 3'b110;
      memory_array[9015] <= 3'b000;
      memory_array[9016] <= 3'b000;
      memory_array[9017] <= 3'b000;
      memory_array[9018] <= 3'b110;
      memory_array[9019] <= 3'b110;
      memory_array[9020] <= 3'b000;
      memory_array[9021] <= 3'b101;
      memory_array[9022] <= 3'b101;
      memory_array[9023] <= 3'b000;
      memory_array[9024] <= 3'b000;
      memory_array[9025] <= 3'b000;
      memory_array[9026] <= 3'b101;
      memory_array[9027] <= 3'b000;
      memory_array[9028] <= 3'b000;
      memory_array[9029] <= 3'b110;
      memory_array[9030] <= 3'b000;
      memory_array[9031] <= 3'b000;
      memory_array[9032] <= 3'b000;
      memory_array[9033] <= 3'b110;
      memory_array[9034] <= 3'b000;
      memory_array[9035] <= 3'b101;
      memory_array[9036] <= 3'b111;
      memory_array[9037] <= 3'b111;
      memory_array[9038] <= 3'b111;
      memory_array[9039] <= 3'b101;
      memory_array[9040] <= 3'b000;
      memory_array[9041] <= 3'b000;
      memory_array[9042] <= 3'b000;
      memory_array[9043] <= 3'b101;
      memory_array[9044] <= 3'b101;
      memory_array[9045] <= 3'b101;
      memory_array[9046] <= 3'b101;
      memory_array[9047] <= 3'b101;
      memory_array[9048] <= 3'b101;
      memory_array[9049] <= 3'b101;
      memory_array[9050] <= 3'b101;
      memory_array[9051] <= 3'b101;
      memory_array[9052] <= 3'b101;
      memory_array[9053] <= 3'b101;
      memory_array[9054] <= 3'b101;
      memory_array[9055] <= 3'b101;
      memory_array[9056] <= 3'b101;
      memory_array[9057] <= 3'b101;
      memory_array[9058] <= 3'b101;
      memory_array[9059] <= 3'b101;
      memory_array[9060] <= 3'b101;
      memory_array[9061] <= 3'b101;
      memory_array[9062] <= 3'b101;
      memory_array[9063] <= 3'b101;
      memory_array[9064] <= 3'b101;
      memory_array[9065] <= 3'b101;
      memory_array[9066] <= 3'b101;
      memory_array[9067] <= 3'b101;
      memory_array[9068] <= 3'b101;
      memory_array[9069] <= 3'b101;
      memory_array[9070] <= 3'b101;
      memory_array[9071] <= 3'b101;
      memory_array[9072] <= 3'b101;
      memory_array[9073] <= 3'b101;
      memory_array[9074] <= 3'b110;
      memory_array[9075] <= 3'b101;
      memory_array[9076] <= 3'b101;
      memory_array[9077] <= 3'b101;
      memory_array[9078] <= 3'b101;
      memory_array[9079] <= 3'b101;
      memory_array[9080] <= 3'b111;
      memory_array[9081] <= 3'b111;
      memory_array[9082] <= 3'b111;
      memory_array[9083] <= 3'b111;
      memory_array[9084] <= 3'b111;
      memory_array[9085] <= 3'b111;
      memory_array[9086] <= 3'b111;
      memory_array[9087] <= 3'b111;
      memory_array[9088] <= 3'b111;
      memory_array[9089] <= 3'b101;
      memory_array[9090] <= 3'b101;
      memory_array[9091] <= 3'b000;
      memory_array[9092] <= 3'b101;
      memory_array[9093] <= 3'b111;
      memory_array[9094] <= 3'b000;
      memory_array[9095] <= 3'b000;
      memory_array[9096] <= 3'b000;
      memory_array[9097] <= 3'b101;
      memory_array[9098] <= 3'b111;
      memory_array[9099] <= 3'b111;
      memory_array[9100] <= 3'b101;
      memory_array[9101] <= 3'b111;
      memory_array[9102] <= 3'b111;
      memory_array[9103] <= 3'b000;
      memory_array[9104] <= 3'b101;
      memory_array[9105] <= 3'b101;
      memory_array[9106] <= 3'b000;
      memory_array[9107] <= 3'b101;
      memory_array[9108] <= 3'b101;
      memory_array[9109] <= 3'b110;
      memory_array[9110] <= 3'b101;
      memory_array[9111] <= 3'b101;
      memory_array[9112] <= 3'b101;
      memory_array[9113] <= 3'b101;
      memory_array[9114] <= 3'b101;
      memory_array[9115] <= 3'b101;
      memory_array[9116] <= 3'b000;
      memory_array[9117] <= 3'b101;
      memory_array[9118] <= 3'b101;
      memory_array[9119] <= 3'b101;
      memory_array[9120] <= 3'b101;
      memory_array[9121] <= 3'b101;
      memory_array[9122] <= 3'b101;
      memory_array[9123] <= 3'b101;
      memory_array[9124] <= 3'b101;
      memory_array[9125] <= 3'b101;
      memory_array[9126] <= 3'b101;
      memory_array[9127] <= 3'b000;
      memory_array[9128] <= 3'b101;
      memory_array[9129] <= 3'b101;
      memory_array[9130] <= 3'b101;
      memory_array[9131] <= 3'b101;
      memory_array[9132] <= 3'b000;
      memory_array[9133] <= 3'b101;
      memory_array[9134] <= 3'b101;
      memory_array[9135] <= 3'b101;
      memory_array[9136] <= 3'b101;
      memory_array[9137] <= 3'b101;
      memory_array[9138] <= 3'b101;
      memory_array[9139] <= 3'b101;
      memory_array[9140] <= 3'b101;
      memory_array[9141] <= 3'b101;
      memory_array[9142] <= 3'b101;
      memory_array[9143] <= 3'b101;
      memory_array[9144] <= 3'b101;
      memory_array[9145] <= 3'b101;
      memory_array[9146] <= 3'b101;
      memory_array[9147] <= 3'b101;
      memory_array[9148] <= 3'b101;
      memory_array[9149] <= 3'b101;
      memory_array[9150] <= 3'b101;
      memory_array[9151] <= 3'b101;
      memory_array[9152] <= 3'b000;
      memory_array[9153] <= 3'b101;
      memory_array[9154] <= 3'b101;
      memory_array[9155] <= 3'b101;
      memory_array[9156] <= 3'b101;
      memory_array[9157] <= 3'b101;
      memory_array[9158] <= 3'b000;
      memory_array[9159] <= 3'b000;
      memory_array[9160] <= 3'b101;
      memory_array[9161] <= 3'b111;
      memory_array[9162] <= 3'b111;
      memory_array[9163] <= 3'b111;
      memory_array[9164] <= 3'b101;
      memory_array[9165] <= 3'b000;
      memory_array[9166] <= 3'b000;
      memory_array[9167] <= 3'b000;
      memory_array[9168] <= 3'b110;
      memory_array[9169] <= 3'b110;
      memory_array[9170] <= 3'b000;
      memory_array[9171] <= 3'b000;
      memory_array[9172] <= 3'b101;
      memory_array[9173] <= 3'b101;
      memory_array[9174] <= 3'b000;
      memory_array[9175] <= 3'b000;
      memory_array[9176] <= 3'b000;
      memory_array[9177] <= 3'b101;
      memory_array[9178] <= 3'b101;
      memory_array[9179] <= 3'b000;
      memory_array[9180] <= 3'b000;
      memory_array[9181] <= 3'b000;
      memory_array[9182] <= 3'b000;
      memory_array[9183] <= 3'b110;
      memory_array[9184] <= 3'b110;
      memory_array[9185] <= 3'b000;
      memory_array[9186] <= 3'b000;
      memory_array[9187] <= 3'b000;
      memory_array[9188] <= 3'b110;
      memory_array[9189] <= 3'b000;
      memory_array[9190] <= 3'b000;
      memory_array[9191] <= 3'b101;
      memory_array[9192] <= 3'b000;
      memory_array[9193] <= 3'b110;
      memory_array[9194] <= 3'b110;
      memory_array[9195] <= 3'b000;
      memory_array[9196] <= 3'b000;
      memory_array[9197] <= 3'b000;
      memory_array[9198] <= 3'b110;
      memory_array[9199] <= 3'b110;
      memory_array[9200] <= 3'b101;
      memory_array[9201] <= 3'b101;
      memory_array[9202] <= 3'b101;
      memory_array[9203] <= 3'b101;
      memory_array[9204] <= 3'b101;
      memory_array[9205] <= 3'b101;
      memory_array[9206] <= 3'b101;
      memory_array[9207] <= 3'b101;
      memory_array[9208] <= 3'b101;
      memory_array[9209] <= 3'b000;
      memory_array[9210] <= 3'b000;
      memory_array[9211] <= 3'b110;
      memory_array[9212] <= 3'b110;
      memory_array[9213] <= 3'b000;
      memory_array[9214] <= 3'b000;
      memory_array[9215] <= 3'b110;
      memory_array[9216] <= 3'b110;
      memory_array[9217] <= 3'b110;
      memory_array[9218] <= 3'b000;
      memory_array[9219] <= 3'b000;
      memory_array[9220] <= 3'b110;
      memory_array[9221] <= 3'b000;
      memory_array[9222] <= 3'b000;
      memory_array[9223] <= 3'b000;
      memory_array[9224] <= 3'b000;
      memory_array[9225] <= 3'b000;
      memory_array[9226] <= 3'b000;
      memory_array[9227] <= 3'b101;
      memory_array[9228] <= 3'b101;
      memory_array[9229] <= 3'b000;
      memory_array[9230] <= 3'b110;
      memory_array[9231] <= 3'b110;
      memory_array[9232] <= 3'b110;
      memory_array[9233] <= 3'b000;
      memory_array[9234] <= 3'b101;
      memory_array[9235] <= 3'b111;
      memory_array[9236] <= 3'b111;
      memory_array[9237] <= 3'b111;
      memory_array[9238] <= 3'b111;
      memory_array[9239] <= 3'b000;
      memory_array[9240] <= 3'b101;
      memory_array[9241] <= 3'b101;
      memory_array[9242] <= 3'b101;
      memory_array[9243] <= 3'b101;
      memory_array[9244] <= 3'b101;
      memory_array[9245] <= 3'b101;
      memory_array[9246] <= 3'b101;
      memory_array[9247] <= 3'b101;
      memory_array[9248] <= 3'b101;
      memory_array[9249] <= 3'b101;
      memory_array[9250] <= 3'b101;
      memory_array[9251] <= 3'b101;
      memory_array[9252] <= 3'b101;
      memory_array[9253] <= 3'b101;
      memory_array[9254] <= 3'b101;
      memory_array[9255] <= 3'b101;
      memory_array[9256] <= 3'b101;
      memory_array[9257] <= 3'b101;
      memory_array[9258] <= 3'b101;
      memory_array[9259] <= 3'b101;
      memory_array[9260] <= 3'b101;
      memory_array[9261] <= 3'b101;
      memory_array[9262] <= 3'b101;
      memory_array[9263] <= 3'b101;
      memory_array[9264] <= 3'b101;
      memory_array[9265] <= 3'b101;
      memory_array[9266] <= 3'b101;
      memory_array[9267] <= 3'b101;
      memory_array[9268] <= 3'b101;
      memory_array[9269] <= 3'b101;
      memory_array[9270] <= 3'b101;
      memory_array[9271] <= 3'b101;
      memory_array[9272] <= 3'b101;
      memory_array[9273] <= 3'b111;
      memory_array[9274] <= 3'b111;
      memory_array[9275] <= 3'b111;
      memory_array[9276] <= 3'b101;
      memory_array[9277] <= 3'b101;
      memory_array[9278] <= 3'b000;
      memory_array[9279] <= 3'b101;
      memory_array[9280] <= 3'b101;
      memory_array[9281] <= 3'b111;
      memory_array[9282] <= 3'b111;
      memory_array[9283] <= 3'b111;
      memory_array[9284] <= 3'b111;
      memory_array[9285] <= 3'b111;
      memory_array[9286] <= 3'b111;
      memory_array[9287] <= 3'b101;
      memory_array[9288] <= 3'b101;
      memory_array[9289] <= 3'b101;
      memory_array[9290] <= 3'b101;
      memory_array[9291] <= 3'b000;
      memory_array[9292] <= 3'b101;
      memory_array[9293] <= 3'b111;
      memory_array[9294] <= 3'b000;
      memory_array[9295] <= 3'b101;
      memory_array[9296] <= 3'b101;
      memory_array[9297] <= 3'b101;
      memory_array[9298] <= 3'b101;
      memory_array[9299] <= 3'b101;
      memory_array[9300] <= 3'b101;
      memory_array[9301] <= 3'b111;
      memory_array[9302] <= 3'b111;
      memory_array[9303] <= 3'b000;
      memory_array[9304] <= 3'b101;
      memory_array[9305] <= 3'b101;
      memory_array[9306] <= 3'b000;
      memory_array[9307] <= 3'b110;
      memory_array[9308] <= 3'b101;
      memory_array[9309] <= 3'b110;
      memory_array[9310] <= 3'b101;
      memory_array[9311] <= 3'b000;
      memory_array[9312] <= 3'b101;
      memory_array[9313] <= 3'b101;
      memory_array[9314] <= 3'b101;
      memory_array[9315] <= 3'b101;
      memory_array[9316] <= 3'b101;
      memory_array[9317] <= 3'b101;
      memory_array[9318] <= 3'b101;
      memory_array[9319] <= 3'b101;
      memory_array[9320] <= 3'b101;
      memory_array[9321] <= 3'b000;
      memory_array[9322] <= 3'b101;
      memory_array[9323] <= 3'b101;
      memory_array[9324] <= 3'b000;
      memory_array[9325] <= 3'b101;
      memory_array[9326] <= 3'b101;
      memory_array[9327] <= 3'b101;
      memory_array[9328] <= 3'b101;
      memory_array[9329] <= 3'b000;
      memory_array[9330] <= 3'b101;
      memory_array[9331] <= 3'b101;
      memory_array[9332] <= 3'b101;
      memory_array[9333] <= 3'b101;
      memory_array[9334] <= 3'b000;
      memory_array[9335] <= 3'b101;
      memory_array[9336] <= 3'b101;
      memory_array[9337] <= 3'b101;
      memory_array[9338] <= 3'b101;
      memory_array[9339] <= 3'b101;
      memory_array[9340] <= 3'b101;
      memory_array[9341] <= 3'b101;
      memory_array[9342] <= 3'b101;
      memory_array[9343] <= 3'b101;
      memory_array[9344] <= 3'b101;
      memory_array[9345] <= 3'b101;
      memory_array[9346] <= 3'b101;
      memory_array[9347] <= 3'b101;
      memory_array[9348] <= 3'b101;
      memory_array[9349] <= 3'b101;
      memory_array[9350] <= 3'b101;
      memory_array[9351] <= 3'b101;
      memory_array[9352] <= 3'b101;
      memory_array[9353] <= 3'b101;
      memory_array[9354] <= 3'b101;
      memory_array[9355] <= 3'b101;
      memory_array[9356] <= 3'b101;
      memory_array[9357] <= 3'b000;
      memory_array[9358] <= 3'b101;
      memory_array[9359] <= 3'b000;
      memory_array[9360] <= 3'b000;
      memory_array[9361] <= 3'b111;
      memory_array[9362] <= 3'b111;
      memory_array[9363] <= 3'b111;
      memory_array[9364] <= 3'b111;
      memory_array[9365] <= 3'b101;
      memory_array[9366] <= 3'b110;
      memory_array[9367] <= 3'b110;
      memory_array[9368] <= 3'b000;
      memory_array[9369] <= 3'b000;
      memory_array[9370] <= 3'b110;
      memory_array[9371] <= 3'b101;
      memory_array[9372] <= 3'b000;
      memory_array[9373] <= 3'b000;
      memory_array[9374] <= 3'b000;
      memory_array[9375] <= 3'b000;
      memory_array[9376] <= 3'b000;
      memory_array[9377] <= 3'b000;
      memory_array[9378] <= 3'b000;
      memory_array[9379] <= 3'b000;
      memory_array[9380] <= 3'b110;
      memory_array[9381] <= 3'b110;
      memory_array[9382] <= 3'b110;
      memory_array[9383] <= 3'b000;
      memory_array[9384] <= 3'b000;
      memory_array[9385] <= 3'b110;
      memory_array[9386] <= 3'b110;
      memory_array[9387] <= 3'b110;
      memory_array[9388] <= 3'b000;
      memory_array[9389] <= 3'b000;
      memory_array[9390] <= 3'b000;
      memory_array[9391] <= 3'b101;
      memory_array[9392] <= 3'b101;
      memory_array[9393] <= 3'b101;
      memory_array[9394] <= 3'b101;
      memory_array[9395] <= 3'b101;
      memory_array[9396] <= 3'b101;
      memory_array[9397] <= 3'b101;
      memory_array[9398] <= 3'b101;
      memory_array[9399] <= 3'b101;
      memory_array[9400] <= 3'b101;
      memory_array[9401] <= 3'b101;
      memory_array[9402] <= 3'b101;
      memory_array[9403] <= 3'b101;
      memory_array[9404] <= 3'b101;
      memory_array[9405] <= 3'b101;
      memory_array[9406] <= 3'b101;
      memory_array[9407] <= 3'b101;
      memory_array[9408] <= 3'b101;
      memory_array[9409] <= 3'b000;
      memory_array[9410] <= 3'b000;
      memory_array[9411] <= 3'b110;
      memory_array[9412] <= 3'b110;
      memory_array[9413] <= 3'b000;
      memory_array[9414] <= 3'b000;
      memory_array[9415] <= 3'b110;
      memory_array[9416] <= 3'b110;
      memory_array[9417] <= 3'b000;
      memory_array[9418] <= 3'b101;
      memory_array[9419] <= 3'b101;
      memory_array[9420] <= 3'b000;
      memory_array[9421] <= 3'b110;
      memory_array[9422] <= 3'b110;
      memory_array[9423] <= 3'b000;
      memory_array[9424] <= 3'b000;
      memory_array[9425] <= 3'b110;
      memory_array[9426] <= 3'b110;
      memory_array[9427] <= 3'b000;
      memory_array[9428] <= 3'b101;
      memory_array[9429] <= 3'b000;
      memory_array[9430] <= 3'b110;
      memory_array[9431] <= 3'b000;
      memory_array[9432] <= 3'b000;
      memory_array[9433] <= 3'b000;
      memory_array[9434] <= 3'b111;
      memory_array[9435] <= 3'b111;
      memory_array[9436] <= 3'b111;
      memory_array[9437] <= 3'b111;
      memory_array[9438] <= 3'b111;
      memory_array[9439] <= 3'b000;
      memory_array[9440] <= 3'b101;
      memory_array[9441] <= 3'b000;
      memory_array[9442] <= 3'b101;
      memory_array[9443] <= 3'b101;
      memory_array[9444] <= 3'b101;
      memory_array[9445] <= 3'b101;
      memory_array[9446] <= 3'b101;
      memory_array[9447] <= 3'b101;
      memory_array[9448] <= 3'b101;
      memory_array[9449] <= 3'b101;
      memory_array[9450] <= 3'b101;
      memory_array[9451] <= 3'b101;
      memory_array[9452] <= 3'b101;
      memory_array[9453] <= 3'b101;
      memory_array[9454] <= 3'b101;
      memory_array[9455] <= 3'b101;
      memory_array[9456] <= 3'b000;
      memory_array[9457] <= 3'b101;
      memory_array[9458] <= 3'b101;
      memory_array[9459] <= 3'b101;
      memory_array[9460] <= 3'b101;
      memory_array[9461] <= 3'b101;
      memory_array[9462] <= 3'b101;
      memory_array[9463] <= 3'b101;
      memory_array[9464] <= 3'b101;
      memory_array[9465] <= 3'b101;
      memory_array[9466] <= 3'b101;
      memory_array[9467] <= 3'b101;
      memory_array[9468] <= 3'b101;
      memory_array[9469] <= 3'b101;
      memory_array[9470] <= 3'b101;
      memory_array[9471] <= 3'b101;
      memory_array[9472] <= 3'b101;
      memory_array[9473] <= 3'b101;
      memory_array[9474] <= 3'b000;
      memory_array[9475] <= 3'b111;
      memory_array[9476] <= 3'b101;
      memory_array[9477] <= 3'b101;
      memory_array[9478] <= 3'b101;
      memory_array[9479] <= 3'b101;
      memory_array[9480] <= 3'b101;
      memory_array[9481] <= 3'b110;
      memory_array[9482] <= 3'b000;
      memory_array[9483] <= 3'b000;
      memory_array[9484] <= 3'b000;
      memory_array[9485] <= 3'b000;
      memory_array[9486] <= 3'b000;
      memory_array[9487] <= 3'b000;
      memory_array[9488] <= 3'b000;
      memory_array[9489] <= 3'b000;
      memory_array[9490] <= 3'b000;
      memory_array[9491] <= 3'b000;
      memory_array[9492] <= 3'b000;
      memory_array[9493] <= 3'b111;
      memory_array[9494] <= 3'b000;
      memory_array[9495] <= 3'b101;
      memory_array[9496] <= 3'b101;
      memory_array[9497] <= 3'b111;
      memory_array[9498] <= 3'b111;
      memory_array[9499] <= 3'b111;
      memory_array[9500] <= 3'b111;
      memory_array[9501] <= 3'b101;
      memory_array[9502] <= 3'b101;
      memory_array[9503] <= 3'b000;
      memory_array[9504] <= 3'b000;
      memory_array[9505] <= 3'b000;
      memory_array[9506] <= 3'b000;
      memory_array[9507] <= 3'b111;
      memory_array[9508] <= 3'b111;
      memory_array[9509] <= 3'b110;
      memory_array[9510] <= 3'b110;
      memory_array[9511] <= 3'b101;
      memory_array[9512] <= 3'b101;
      memory_array[9513] <= 3'b101;
      memory_array[9514] <= 3'b101;
      memory_array[9515] <= 3'b101;
      memory_array[9516] <= 3'b101;
      memory_array[9517] <= 3'b101;
      memory_array[9518] <= 3'b101;
      memory_array[9519] <= 3'b101;
      memory_array[9520] <= 3'b101;
      memory_array[9521] <= 3'b101;
      memory_array[9522] <= 3'b101;
      memory_array[9523] <= 3'b101;
      memory_array[9524] <= 3'b101;
      memory_array[9525] <= 3'b101;
      memory_array[9526] <= 3'b101;
      memory_array[9527] <= 3'b101;
      memory_array[9528] <= 3'b101;
      memory_array[9529] <= 3'b101;
      memory_array[9530] <= 3'b101;
      memory_array[9531] <= 3'b101;
      memory_array[9532] <= 3'b101;
      memory_array[9533] <= 3'b101;
      memory_array[9534] <= 3'b000;
      memory_array[9535] <= 3'b000;
      memory_array[9536] <= 3'b101;
      memory_array[9537] <= 3'b101;
      memory_array[9538] <= 3'b101;
      memory_array[9539] <= 3'b101;
      memory_array[9540] <= 3'b101;
      memory_array[9541] <= 3'b101;
      memory_array[9542] <= 3'b101;
      memory_array[9543] <= 3'b000;
      memory_array[9544] <= 3'b101;
      memory_array[9545] <= 3'b101;
      memory_array[9546] <= 3'b110;
      memory_array[9547] <= 3'b101;
      memory_array[9548] <= 3'b101;
      memory_array[9549] <= 3'b101;
      memory_array[9550] <= 3'b101;
      memory_array[9551] <= 3'b101;
      memory_array[9552] <= 3'b101;
      memory_array[9553] <= 3'b101;
      memory_array[9554] <= 3'b101;
      memory_array[9555] <= 3'b101;
      memory_array[9556] <= 3'b101;
      memory_array[9557] <= 3'b101;
      memory_array[9558] <= 3'b000;
      memory_array[9559] <= 3'b101;
      memory_array[9560] <= 3'b000;
      memory_array[9561] <= 3'b111;
      memory_array[9562] <= 3'b111;
      memory_array[9563] <= 3'b111;
      memory_array[9564] <= 3'b111;
      memory_array[9565] <= 3'b111;
      memory_array[9566] <= 3'b000;
      memory_array[9567] <= 3'b101;
      memory_array[9568] <= 3'b000;
      memory_array[9569] <= 3'b000;
      memory_array[9570] <= 3'b110;
      memory_array[9571] <= 3'b101;
      memory_array[9572] <= 3'b000;
      memory_array[9573] <= 3'b000;
      memory_array[9574] <= 3'b000;
      memory_array[9575] <= 3'b110;
      memory_array[9576] <= 3'b110;
      memory_array[9577] <= 3'b110;
      memory_array[9578] <= 3'b000;
      memory_array[9579] <= 3'b000;
      memory_array[9580] <= 3'b101;
      memory_array[9581] <= 3'b101;
      memory_array[9582] <= 3'b110;
      memory_array[9583] <= 3'b000;
      memory_array[9584] <= 3'b000;
      memory_array[9585] <= 3'b110;
      memory_array[9586] <= 3'b110;
      memory_array[9587] <= 3'b110;
      memory_array[9588] <= 3'b000;
      memory_array[9589] <= 3'b000;
      memory_array[9590] <= 3'b000;
      memory_array[9591] <= 3'b101;
      memory_array[9592] <= 3'b101;
      memory_array[9593] <= 3'b101;
      memory_array[9594] <= 3'b101;
      memory_array[9595] <= 3'b101;
      memory_array[9596] <= 3'b101;
      memory_array[9597] <= 3'b101;
      memory_array[9598] <= 3'b101;
      memory_array[9599] <= 3'b101;
      memory_array[9600] <= 3'b000;
      memory_array[9601] <= 3'b000;
      memory_array[9602] <= 3'b000;
      memory_array[9603] <= 3'b110;
      memory_array[9604] <= 3'b110;
      memory_array[9605] <= 3'b000;
      memory_array[9606] <= 3'b000;
      memory_array[9607] <= 3'b000;
      memory_array[9608] <= 3'b101;
      memory_array[9609] <= 3'b000;
      memory_array[9610] <= 3'b000;
      memory_array[9611] <= 3'b000;
      memory_array[9612] <= 3'b000;
      memory_array[9613] <= 3'b110;
      memory_array[9614] <= 3'b101;
      memory_array[9615] <= 3'b101;
      memory_array[9616] <= 3'b000;
      memory_array[9617] <= 3'b101;
      memory_array[9618] <= 3'b101;
      memory_array[9619] <= 3'b101;
      memory_array[9620] <= 3'b101;
      memory_array[9621] <= 3'b000;
      memory_array[9622] <= 3'b000;
      memory_array[9623] <= 3'b110;
      memory_array[9624] <= 3'b110;
      memory_array[9625] <= 3'b000;
      memory_array[9626] <= 3'b000;
      memory_array[9627] <= 3'b101;
      memory_array[9628] <= 3'b101;
      memory_array[9629] <= 3'b000;
      memory_array[9630] <= 3'b000;
      memory_array[9631] <= 3'b000;
      memory_array[9632] <= 3'b101;
      memory_array[9633] <= 3'b000;
      memory_array[9634] <= 3'b111;
      memory_array[9635] <= 3'b111;
      memory_array[9636] <= 3'b111;
      memory_array[9637] <= 3'b111;
      memory_array[9638] <= 3'b111;
      memory_array[9639] <= 3'b101;
      memory_array[9640] <= 3'b101;
      memory_array[9641] <= 3'b000;
      memory_array[9642] <= 3'b101;
      memory_array[9643] <= 3'b101;
      memory_array[9644] <= 3'b101;
      memory_array[9645] <= 3'b101;
      memory_array[9646] <= 3'b101;
      memory_array[9647] <= 3'b101;
      memory_array[9648] <= 3'b101;
      memory_array[9649] <= 3'b101;
      memory_array[9650] <= 3'b101;
      memory_array[9651] <= 3'b101;
      memory_array[9652] <= 3'b101;
      memory_array[9653] <= 3'b101;
      memory_array[9654] <= 3'b101;
      memory_array[9655] <= 3'b101;
      memory_array[9656] <= 3'b101;
      memory_array[9657] <= 3'b101;
      memory_array[9658] <= 3'b101;
      memory_array[9659] <= 3'b101;
      memory_array[9660] <= 3'b101;
      memory_array[9661] <= 3'b101;
      memory_array[9662] <= 3'b101;
      memory_array[9663] <= 3'b101;
      memory_array[9664] <= 3'b101;
      memory_array[9665] <= 3'b101;
      memory_array[9666] <= 3'b101;
      memory_array[9667] <= 3'b101;
      memory_array[9668] <= 3'b101;
      memory_array[9669] <= 3'b101;
      memory_array[9670] <= 3'b101;
      memory_array[9671] <= 3'b101;
      memory_array[9672] <= 3'b101;
      memory_array[9673] <= 3'b101;
      memory_array[9674] <= 3'b000;
      memory_array[9675] <= 3'b111;
      memory_array[9676] <= 3'b101;
      memory_array[9677] <= 3'b101;
      memory_array[9678] <= 3'b101;
      memory_array[9679] <= 3'b101;
      memory_array[9680] <= 3'b101;
      memory_array[9681] <= 3'b101;
      memory_array[9682] <= 3'b000;
      memory_array[9683] <= 3'b111;
      memory_array[9684] <= 3'b111;
      memory_array[9685] <= 3'b000;
      memory_array[9686] <= 3'b000;
      memory_array[9687] <= 3'b000;
      memory_array[9688] <= 3'b111;
      memory_array[9689] <= 3'b000;
      memory_array[9690] <= 3'b000;
      memory_array[9691] <= 3'b000;
      memory_array[9692] <= 3'b000;
      memory_array[9693] <= 3'b111;
      memory_array[9694] <= 3'b000;
      memory_array[9695] <= 3'b000;
      memory_array[9696] <= 3'b000;
      memory_array[9697] <= 3'b101;
      memory_array[9698] <= 3'b111;
      memory_array[9699] <= 3'b111;
      memory_array[9700] <= 3'b111;
      memory_array[9701] <= 3'b111;
      memory_array[9702] <= 3'b111;
      memory_array[9703] <= 3'b101;
      memory_array[9704] <= 3'b101;
      memory_array[9705] <= 3'b000;
      memory_array[9706] <= 3'b000;
      memory_array[9707] <= 3'b111;
      memory_array[9708] <= 3'b110;
      memory_array[9709] <= 3'b000;
      memory_array[9710] <= 3'b101;
      memory_array[9711] <= 3'b110;
      memory_array[9712] <= 3'b101;
      memory_array[9713] <= 3'b101;
      memory_array[9714] <= 3'b101;
      memory_array[9715] <= 3'b101;
      memory_array[9716] <= 3'b101;
      memory_array[9717] <= 3'b101;
      memory_array[9718] <= 3'b101;
      memory_array[9719] <= 3'b101;
      memory_array[9720] <= 3'b101;
      memory_array[9721] <= 3'b101;
      memory_array[9722] <= 3'b101;
      memory_array[9723] <= 3'b101;
      memory_array[9724] <= 3'b101;
      memory_array[9725] <= 3'b101;
      memory_array[9726] <= 3'b101;
      memory_array[9727] <= 3'b101;
      memory_array[9728] <= 3'b101;
      memory_array[9729] <= 3'b101;
      memory_array[9730] <= 3'b101;
      memory_array[9731] <= 3'b101;
      memory_array[9732] <= 3'b101;
      memory_array[9733] <= 3'b101;
      memory_array[9734] <= 3'b101;
      memory_array[9735] <= 3'b101;
      memory_array[9736] <= 3'b101;
      memory_array[9737] <= 3'b101;
      memory_array[9738] <= 3'b101;
      memory_array[9739] <= 3'b101;
      memory_array[9740] <= 3'b101;
      memory_array[9741] <= 3'b101;
      memory_array[9742] <= 3'b000;
      memory_array[9743] <= 3'b101;
      memory_array[9744] <= 3'b101;
      memory_array[9745] <= 3'b110;
      memory_array[9746] <= 3'b101;
      memory_array[9747] <= 3'b101;
      memory_array[9748] <= 3'b101;
      memory_array[9749] <= 3'b101;
      memory_array[9750] <= 3'b101;
      memory_array[9751] <= 3'b101;
      memory_array[9752] <= 3'b101;
      memory_array[9753] <= 3'b101;
      memory_array[9754] <= 3'b101;
      memory_array[9755] <= 3'b101;
      memory_array[9756] <= 3'b101;
      memory_array[9757] <= 3'b101;
      memory_array[9758] <= 3'b000;
      memory_array[9759] <= 3'b101;
      memory_array[9760] <= 3'b000;
      memory_array[9761] <= 3'b111;
      memory_array[9762] <= 3'b111;
      memory_array[9763] <= 3'b111;
      memory_array[9764] <= 3'b111;
      memory_array[9765] <= 3'b111;
      memory_array[9766] <= 3'b000;
      memory_array[9767] <= 3'b000;
      memory_array[9768] <= 3'b000;
      memory_array[9769] <= 3'b000;
      memory_array[9770] <= 3'b000;
      memory_array[9771] <= 3'b101;
      memory_array[9772] <= 3'b000;
      memory_array[9773] <= 3'b110;
      memory_array[9774] <= 3'b110;
      memory_array[9775] <= 3'b000;
      memory_array[9776] <= 3'b000;
      memory_array[9777] <= 3'b000;
      memory_array[9778] <= 3'b110;
      memory_array[9779] <= 3'b101;
      memory_array[9780] <= 3'b101;
      memory_array[9781] <= 3'b101;
      memory_array[9782] <= 3'b000;
      memory_array[9783] <= 3'b110;
      memory_array[9784] <= 3'b101;
      memory_array[9785] <= 3'b101;
      memory_array[9786] <= 3'b000;
      memory_array[9787] <= 3'b000;
      memory_array[9788] <= 3'b110;
      memory_array[9789] <= 3'b000;
      memory_array[9790] <= 3'b000;
      memory_array[9791] <= 3'b101;
      memory_array[9792] <= 3'b000;
      memory_array[9793] <= 3'b110;
      memory_array[9794] <= 3'b110;
      memory_array[9795] <= 3'b000;
      memory_array[9796] <= 3'b000;
      memory_array[9797] <= 3'b000;
      memory_array[9798] <= 3'b110;
      memory_array[9799] <= 3'b110;
      memory_array[9800] <= 3'b101;
      memory_array[9801] <= 3'b000;
      memory_array[9802] <= 3'b000;
      memory_array[9803] <= 3'b110;
      memory_array[9804] <= 3'b110;
      memory_array[9805] <= 3'b000;
      memory_array[9806] <= 3'b101;
      memory_array[9807] <= 3'b101;
      memory_array[9808] <= 3'b101;
      memory_array[9809] <= 3'b000;
      memory_array[9810] <= 3'b000;
      memory_array[9811] <= 3'b000;
      memory_array[9812] <= 3'b000;
      memory_array[9813] <= 3'b000;
      memory_array[9814] <= 3'b000;
      memory_array[9815] <= 3'b000;
      memory_array[9816] <= 3'b000;
      memory_array[9817] <= 3'b101;
      memory_array[9818] <= 3'b101;
      memory_array[9819] <= 3'b101;
      memory_array[9820] <= 3'b101;
      memory_array[9821] <= 3'b000;
      memory_array[9822] <= 3'b000;
      memory_array[9823] <= 3'b110;
      memory_array[9824] <= 3'b110;
      memory_array[9825] <= 3'b000;
      memory_array[9826] <= 3'b000;
      memory_array[9827] <= 3'b000;
      memory_array[9828] <= 3'b000;
      memory_array[9829] <= 3'b101;
      memory_array[9830] <= 3'b000;
      memory_array[9831] <= 3'b000;
      memory_array[9832] <= 3'b101;
      memory_array[9833] <= 3'b000;
      memory_array[9834] <= 3'b111;
      memory_array[9835] <= 3'b111;
      memory_array[9836] <= 3'b111;
      memory_array[9837] <= 3'b111;
      memory_array[9838] <= 3'b101;
      memory_array[9839] <= 3'b101;
      memory_array[9840] <= 3'b101;
      memory_array[9841] <= 3'b101;
      memory_array[9842] <= 3'b101;
      memory_array[9843] <= 3'b101;
      memory_array[9844] <= 3'b101;
      memory_array[9845] <= 3'b101;
      memory_array[9846] <= 3'b101;
      memory_array[9847] <= 3'b101;
      memory_array[9848] <= 3'b101;
      memory_array[9849] <= 3'b101;
      memory_array[9850] <= 3'b101;
      memory_array[9851] <= 3'b101;
      memory_array[9852] <= 3'b101;
      memory_array[9853] <= 3'b101;
      memory_array[9854] <= 3'b101;
      memory_array[9855] <= 3'b101;
      memory_array[9856] <= 3'b101;
      memory_array[9857] <= 3'b101;
      memory_array[9858] <= 3'b101;
      memory_array[9859] <= 3'b101;
      memory_array[9860] <= 3'b101;
      memory_array[9861] <= 3'b101;
      memory_array[9862] <= 3'b101;
      memory_array[9863] <= 3'b101;
      memory_array[9864] <= 3'b101;
      memory_array[9865] <= 3'b101;
      memory_array[9866] <= 3'b101;
      memory_array[9867] <= 3'b101;
      memory_array[9868] <= 3'b101;
      memory_array[9869] <= 3'b101;
      memory_array[9870] <= 3'b101;
      memory_array[9871] <= 3'b101;
      memory_array[9872] <= 3'b101;
      memory_array[9873] <= 3'b101;
      memory_array[9874] <= 3'b101;
      memory_array[9875] <= 3'b111;
      memory_array[9876] <= 3'b101;
      memory_array[9877] <= 3'b101;
      memory_array[9878] <= 3'b101;
      memory_array[9879] <= 3'b101;
      memory_array[9880] <= 3'b101;
      memory_array[9881] <= 3'b111;
      memory_array[9882] <= 3'b111;
      memory_array[9883] <= 3'b111;
      memory_array[9884] <= 3'b111;
      memory_array[9885] <= 3'b111;
      memory_array[9886] <= 3'b111;
      memory_array[9887] <= 3'b111;
      memory_array[9888] <= 3'b111;
      memory_array[9889] <= 3'b000;
      memory_array[9890] <= 3'b000;
      memory_array[9891] <= 3'b000;
      memory_array[9892] <= 3'b000;
      memory_array[9893] <= 3'b000;
      memory_array[9894] <= 3'b000;
      memory_array[9895] <= 3'b000;
      memory_array[9896] <= 3'b000;
      memory_array[9897] <= 3'b000;
      memory_array[9898] <= 3'b101;
      memory_array[9899] <= 3'b101;
      memory_array[9900] <= 3'b101;
      memory_array[9901] <= 3'b101;
      memory_array[9902] <= 3'b111;
      memory_array[9903] <= 3'b111;
      memory_array[9904] <= 3'b101;
      memory_array[9905] <= 3'b101;
      memory_array[9906] <= 3'b101;
      memory_array[9907] <= 3'b101;
      memory_array[9908] <= 3'b101;
      memory_array[9909] <= 3'b000;
      memory_array[9910] <= 3'b000;
      memory_array[9911] <= 3'b101;
      memory_array[9912] <= 3'b101;
      memory_array[9913] <= 3'b101;
      memory_array[9914] <= 3'b101;
      memory_array[9915] <= 3'b101;
      memory_array[9916] <= 3'b101;
      memory_array[9917] <= 3'b101;
      memory_array[9918] <= 3'b111;
      memory_array[9919] <= 3'b111;
      memory_array[9920] <= 3'b000;
      memory_array[9921] <= 3'b101;
      memory_array[9922] <= 3'b101;
      memory_array[9923] <= 3'b101;
      memory_array[9924] <= 3'b101;
      memory_array[9925] <= 3'b101;
      memory_array[9926] <= 3'b101;
      memory_array[9927] <= 3'b101;
      memory_array[9928] <= 3'b101;
      memory_array[9929] <= 3'b000;
      memory_array[9930] <= 3'b101;
      memory_array[9931] <= 3'b101;
      memory_array[9932] <= 3'b101;
      memory_array[9933] <= 3'b101;
      memory_array[9934] <= 3'b101;
      memory_array[9935] <= 3'b101;
      memory_array[9936] <= 3'b101;
      memory_array[9937] <= 3'b101;
      memory_array[9938] <= 3'b101;
      memory_array[9939] <= 3'b101;
      memory_array[9940] <= 3'b101;
      memory_array[9941] <= 3'b101;
      memory_array[9942] <= 3'b110;
      memory_array[9943] <= 3'b101;
      memory_array[9944] <= 3'b110;
      memory_array[9945] <= 3'b110;
      memory_array[9946] <= 3'b110;
      memory_array[9947] <= 3'b000;
      memory_array[9948] <= 3'b110;
      memory_array[9949] <= 3'b101;
      memory_array[9950] <= 3'b101;
      memory_array[9951] <= 3'b101;
      memory_array[9952] <= 3'b101;
      memory_array[9953] <= 3'b101;
      memory_array[9954] <= 3'b101;
      memory_array[9955] <= 3'b101;
      memory_array[9956] <= 3'b101;
      memory_array[9957] <= 3'b101;
      memory_array[9958] <= 3'b101;
      memory_array[9959] <= 3'b101;
      memory_array[9960] <= 3'b101;
      memory_array[9961] <= 3'b101;
      memory_array[9962] <= 3'b111;
      memory_array[9963] <= 3'b111;
      memory_array[9964] <= 3'b111;
      memory_array[9965] <= 3'b111;
      memory_array[9966] <= 3'b000;
      memory_array[9967] <= 3'b000;
      memory_array[9968] <= 3'b110;
      memory_array[9969] <= 3'b000;
      memory_array[9970] <= 3'b101;
      memory_array[9971] <= 3'b000;
      memory_array[9972] <= 3'b000;
      memory_array[9973] <= 3'b110;
      memory_array[9974] <= 3'b110;
      memory_array[9975] <= 3'b000;
      memory_array[9976] <= 3'b000;
      memory_array[9977] <= 3'b000;
      memory_array[9978] <= 3'b110;
      memory_array[9979] <= 3'b101;
      memory_array[9980] <= 3'b101;
      memory_array[9981] <= 3'b101;
      memory_array[9982] <= 3'b000;
      memory_array[9983] <= 3'b000;
      memory_array[9984] <= 3'b000;
      memory_array[9985] <= 3'b000;
      memory_array[9986] <= 3'b000;
      memory_array[9987] <= 3'b000;
      memory_array[9988] <= 3'b110;
      memory_array[9989] <= 3'b000;
      memory_array[9990] <= 3'b000;
      memory_array[9991] <= 3'b101;
      memory_array[9992] <= 3'b101;
      memory_array[9993] <= 3'b110;
      memory_array[9994] <= 3'b110;
      memory_array[9995] <= 3'b000;
      memory_array[9996] <= 3'b000;
      memory_array[9997] <= 3'b000;
      memory_array[9998] <= 3'b110;
      memory_array[9999] <= 3'b101;
      memory_array[10000] <= 3'b101;
      memory_array[10001] <= 3'b000;
      memory_array[10002] <= 3'b000;
      memory_array[10003] <= 3'b110;
      memory_array[10004] <= 3'b110;
      memory_array[10005] <= 3'b000;
      memory_array[10006] <= 3'b101;
      memory_array[10007] <= 3'b101;
      memory_array[10008] <= 3'b101;
      memory_array[10009] <= 3'b000;
      memory_array[10010] <= 3'b000;
      memory_array[10011] <= 3'b000;
      memory_array[10012] <= 3'b000;
      memory_array[10013] <= 3'b000;
      memory_array[10014] <= 3'b000;
      memory_array[10015] <= 3'b000;
      memory_array[10016] <= 3'b000;
      memory_array[10017] <= 3'b101;
      memory_array[10018] <= 3'b101;
      memory_array[10019] <= 3'b101;
      memory_array[10020] <= 3'b101;
      memory_array[10021] <= 3'b000;
      memory_array[10022] <= 3'b000;
      memory_array[10023] <= 3'b110;
      memory_array[10024] <= 3'b110;
      memory_array[10025] <= 3'b000;
      memory_array[10026] <= 3'b000;
      memory_array[10027] <= 3'b000;
      memory_array[10028] <= 3'b000;
      memory_array[10029] <= 3'b101;
      memory_array[10030] <= 3'b000;
      memory_array[10031] <= 3'b000;
      memory_array[10032] <= 3'b101;
      memory_array[10033] <= 3'b000;
      memory_array[10034] <= 3'b111;
      memory_array[10035] <= 3'b111;
      memory_array[10036] <= 3'b111;
      memory_array[10037] <= 3'b111;
      memory_array[10038] <= 3'b101;
      memory_array[10039] <= 3'b101;
      memory_array[10040] <= 3'b101;
      memory_array[10041] <= 3'b101;
      memory_array[10042] <= 3'b101;
      memory_array[10043] <= 3'b101;
      memory_array[10044] <= 3'b101;
      memory_array[10045] <= 3'b101;
      memory_array[10046] <= 3'b101;
      memory_array[10047] <= 3'b101;
      memory_array[10048] <= 3'b101;
      memory_array[10049] <= 3'b101;
      memory_array[10050] <= 3'b101;
      memory_array[10051] <= 3'b101;
      memory_array[10052] <= 3'b101;
      memory_array[10053] <= 3'b101;
      memory_array[10054] <= 3'b101;
      memory_array[10055] <= 3'b101;
      memory_array[10056] <= 3'b101;
      memory_array[10057] <= 3'b101;
      memory_array[10058] <= 3'b101;
      memory_array[10059] <= 3'b101;
      memory_array[10060] <= 3'b101;
      memory_array[10061] <= 3'b101;
      memory_array[10062] <= 3'b101;
      memory_array[10063] <= 3'b101;
      memory_array[10064] <= 3'b101;
      memory_array[10065] <= 3'b101;
      memory_array[10066] <= 3'b101;
      memory_array[10067] <= 3'b101;
      memory_array[10068] <= 3'b101;
      memory_array[10069] <= 3'b101;
      memory_array[10070] <= 3'b101;
      memory_array[10071] <= 3'b101;
      memory_array[10072] <= 3'b101;
      memory_array[10073] <= 3'b101;
      memory_array[10074] <= 3'b101;
      memory_array[10075] <= 3'b111;
      memory_array[10076] <= 3'b101;
      memory_array[10077] <= 3'b101;
      memory_array[10078] <= 3'b101;
      memory_array[10079] <= 3'b101;
      memory_array[10080] <= 3'b101;
      memory_array[10081] <= 3'b111;
      memory_array[10082] <= 3'b111;
      memory_array[10083] <= 3'b111;
      memory_array[10084] <= 3'b111;
      memory_array[10085] <= 3'b111;
      memory_array[10086] <= 3'b111;
      memory_array[10087] <= 3'b111;
      memory_array[10088] <= 3'b111;
      memory_array[10089] <= 3'b000;
      memory_array[10090] <= 3'b000;
      memory_array[10091] <= 3'b000;
      memory_array[10092] <= 3'b000;
      memory_array[10093] <= 3'b000;
      memory_array[10094] <= 3'b000;
      memory_array[10095] <= 3'b000;
      memory_array[10096] <= 3'b000;
      memory_array[10097] <= 3'b000;
      memory_array[10098] <= 3'b101;
      memory_array[10099] <= 3'b101;
      memory_array[10100] <= 3'b101;
      memory_array[10101] <= 3'b101;
      memory_array[10102] <= 3'b111;
      memory_array[10103] <= 3'b111;
      memory_array[10104] <= 3'b101;
      memory_array[10105] <= 3'b101;
      memory_array[10106] <= 3'b101;
      memory_array[10107] <= 3'b101;
      memory_array[10108] <= 3'b101;
      memory_array[10109] <= 3'b000;
      memory_array[10110] <= 3'b000;
      memory_array[10111] <= 3'b101;
      memory_array[10112] <= 3'b101;
      memory_array[10113] <= 3'b101;
      memory_array[10114] <= 3'b101;
      memory_array[10115] <= 3'b101;
      memory_array[10116] <= 3'b101;
      memory_array[10117] <= 3'b101;
      memory_array[10118] <= 3'b111;
      memory_array[10119] <= 3'b111;
      memory_array[10120] <= 3'b000;
      memory_array[10121] <= 3'b101;
      memory_array[10122] <= 3'b101;
      memory_array[10123] <= 3'b101;
      memory_array[10124] <= 3'b101;
      memory_array[10125] <= 3'b101;
      memory_array[10126] <= 3'b101;
      memory_array[10127] <= 3'b101;
      memory_array[10128] <= 3'b101;
      memory_array[10129] <= 3'b000;
      memory_array[10130] <= 3'b101;
      memory_array[10131] <= 3'b101;
      memory_array[10132] <= 3'b101;
      memory_array[10133] <= 3'b101;
      memory_array[10134] <= 3'b101;
      memory_array[10135] <= 3'b101;
      memory_array[10136] <= 3'b101;
      memory_array[10137] <= 3'b101;
      memory_array[10138] <= 3'b101;
      memory_array[10139] <= 3'b101;
      memory_array[10140] <= 3'b101;
      memory_array[10141] <= 3'b101;
      memory_array[10142] <= 3'b110;
      memory_array[10143] <= 3'b101;
      memory_array[10144] <= 3'b110;
      memory_array[10145] <= 3'b110;
      memory_array[10146] <= 3'b110;
      memory_array[10147] <= 3'b000;
      memory_array[10148] <= 3'b110;
      memory_array[10149] <= 3'b101;
      memory_array[10150] <= 3'b101;
      memory_array[10151] <= 3'b101;
      memory_array[10152] <= 3'b101;
      memory_array[10153] <= 3'b101;
      memory_array[10154] <= 3'b101;
      memory_array[10155] <= 3'b101;
      memory_array[10156] <= 3'b101;
      memory_array[10157] <= 3'b101;
      memory_array[10158] <= 3'b101;
      memory_array[10159] <= 3'b101;
      memory_array[10160] <= 3'b101;
      memory_array[10161] <= 3'b101;
      memory_array[10162] <= 3'b111;
      memory_array[10163] <= 3'b111;
      memory_array[10164] <= 3'b111;
      memory_array[10165] <= 3'b111;
      memory_array[10166] <= 3'b000;
      memory_array[10167] <= 3'b000;
      memory_array[10168] <= 3'b110;
      memory_array[10169] <= 3'b000;
      memory_array[10170] <= 3'b101;
      memory_array[10171] <= 3'b000;
      memory_array[10172] <= 3'b000;
      memory_array[10173] <= 3'b110;
      memory_array[10174] <= 3'b110;
      memory_array[10175] <= 3'b000;
      memory_array[10176] <= 3'b000;
      memory_array[10177] <= 3'b000;
      memory_array[10178] <= 3'b110;
      memory_array[10179] <= 3'b101;
      memory_array[10180] <= 3'b101;
      memory_array[10181] <= 3'b101;
      memory_array[10182] <= 3'b000;
      memory_array[10183] <= 3'b000;
      memory_array[10184] <= 3'b000;
      memory_array[10185] <= 3'b000;
      memory_array[10186] <= 3'b000;
      memory_array[10187] <= 3'b000;
      memory_array[10188] <= 3'b110;
      memory_array[10189] <= 3'b000;
      memory_array[10190] <= 3'b000;
      memory_array[10191] <= 3'b101;
      memory_array[10192] <= 3'b101;
      memory_array[10193] <= 3'b110;
      memory_array[10194] <= 3'b110;
      memory_array[10195] <= 3'b000;
      memory_array[10196] <= 3'b000;
      memory_array[10197] <= 3'b000;
      memory_array[10198] <= 3'b110;
      memory_array[10199] <= 3'b101;
      memory_array[10200] <= 3'b101;
      memory_array[10201] <= 3'b101;
      memory_array[10202] <= 3'b101;
      memory_array[10203] <= 3'b111;
      memory_array[10204] <= 3'b111;
      memory_array[10205] <= 3'b101;
      memory_array[10206] <= 3'b101;
      memory_array[10207] <= 3'b101;
      memory_array[10208] <= 3'b101;
      memory_array[10209] <= 3'b000;
      memory_array[10210] <= 3'b000;
      memory_array[10211] <= 3'b000;
      memory_array[10212] <= 3'b000;
      memory_array[10213] <= 3'b101;
      memory_array[10214] <= 3'b110;
      memory_array[10215] <= 3'b000;
      memory_array[10216] <= 3'b000;
      memory_array[10217] <= 3'b000;
      memory_array[10218] <= 3'b000;
      memory_array[10219] <= 3'b000;
      memory_array[10220] <= 3'b000;
      memory_array[10221] <= 3'b000;
      memory_array[10222] <= 3'b000;
      memory_array[10223] <= 3'b110;
      memory_array[10224] <= 3'b110;
      memory_array[10225] <= 3'b000;
      memory_array[10226] <= 3'b101;
      memory_array[10227] <= 3'b000;
      memory_array[10228] <= 3'b110;
      memory_array[10229] <= 3'b110;
      memory_array[10230] <= 3'b000;
      memory_array[10231] <= 3'b000;
      memory_array[10232] <= 3'b000;
      memory_array[10233] <= 3'b000;
      memory_array[10234] <= 3'b111;
      memory_array[10235] <= 3'b111;
      memory_array[10236] <= 3'b111;
      memory_array[10237] <= 3'b111;
      memory_array[10238] <= 3'b000;
      memory_array[10239] <= 3'b101;
      memory_array[10240] <= 3'b101;
      memory_array[10241] <= 3'b101;
      memory_array[10242] <= 3'b101;
      memory_array[10243] <= 3'b101;
      memory_array[10244] <= 3'b101;
      memory_array[10245] <= 3'b101;
      memory_array[10246] <= 3'b101;
      memory_array[10247] <= 3'b101;
      memory_array[10248] <= 3'b101;
      memory_array[10249] <= 3'b101;
      memory_array[10250] <= 3'b101;
      memory_array[10251] <= 3'b101;
      memory_array[10252] <= 3'b101;
      memory_array[10253] <= 3'b101;
      memory_array[10254] <= 3'b101;
      memory_array[10255] <= 3'b101;
      memory_array[10256] <= 3'b101;
      memory_array[10257] <= 3'b101;
      memory_array[10258] <= 3'b101;
      memory_array[10259] <= 3'b101;
      memory_array[10260] <= 3'b101;
      memory_array[10261] <= 3'b101;
      memory_array[10262] <= 3'b101;
      memory_array[10263] <= 3'b101;
      memory_array[10264] <= 3'b101;
      memory_array[10265] <= 3'b101;
      memory_array[10266] <= 3'b101;
      memory_array[10267] <= 3'b101;
      memory_array[10268] <= 3'b101;
      memory_array[10269] <= 3'b101;
      memory_array[10270] <= 3'b101;
      memory_array[10271] <= 3'b101;
      memory_array[10272] <= 3'b101;
      memory_array[10273] <= 3'b101;
      memory_array[10274] <= 3'b110;
      memory_array[10275] <= 3'b110;
      memory_array[10276] <= 3'b000;
      memory_array[10277] <= 3'b101;
      memory_array[10278] <= 3'b101;
      memory_array[10279] <= 3'b101;
      memory_array[10280] <= 3'b000;
      memory_array[10281] <= 3'b111;
      memory_array[10282] <= 3'b111;
      memory_array[10283] <= 3'b111;
      memory_array[10284] <= 3'b111;
      memory_array[10285] <= 3'b111;
      memory_array[10286] <= 3'b111;
      memory_array[10287] <= 3'b111;
      memory_array[10288] <= 3'b111;
      memory_array[10289] <= 3'b111;
      memory_array[10290] <= 3'b101;
      memory_array[10291] <= 3'b000;
      memory_array[10292] <= 3'b000;
      memory_array[10293] <= 3'b000;
      memory_array[10294] <= 3'b000;
      memory_array[10295] <= 3'b000;
      memory_array[10296] <= 3'b000;
      memory_array[10297] <= 3'b000;
      memory_array[10298] <= 3'b110;
      memory_array[10299] <= 3'b110;
      memory_array[10300] <= 3'b000;
      memory_array[10301] <= 3'b101;
      memory_array[10302] <= 3'b101;
      memory_array[10303] <= 3'b110;
      memory_array[10304] <= 3'b101;
      memory_array[10305] <= 3'b101;
      memory_array[10306] <= 3'b111;
      memory_array[10307] <= 3'b111;
      memory_array[10308] <= 3'b111;
      memory_array[10309] <= 3'b101;
      memory_array[10310] <= 3'b000;
      memory_array[10311] <= 3'b101;
      memory_array[10312] <= 3'b101;
      memory_array[10313] <= 3'b101;
      memory_array[10314] <= 3'b101;
      memory_array[10315] <= 3'b101;
      memory_array[10316] <= 3'b101;
      memory_array[10317] <= 3'b101;
      memory_array[10318] <= 3'b101;
      memory_array[10319] <= 3'b101;
      memory_array[10320] <= 3'b101;
      memory_array[10321] <= 3'b101;
      memory_array[10322] <= 3'b101;
      memory_array[10323] <= 3'b101;
      memory_array[10324] <= 3'b101;
      memory_array[10325] <= 3'b101;
      memory_array[10326] <= 3'b101;
      memory_array[10327] <= 3'b101;
      memory_array[10328] <= 3'b101;
      memory_array[10329] <= 3'b101;
      memory_array[10330] <= 3'b101;
      memory_array[10331] <= 3'b101;
      memory_array[10332] <= 3'b110;
      memory_array[10333] <= 3'b101;
      memory_array[10334] <= 3'b101;
      memory_array[10335] <= 3'b101;
      memory_array[10336] <= 3'b101;
      memory_array[10337] <= 3'b101;
      memory_array[10338] <= 3'b101;
      memory_array[10339] <= 3'b101;
      memory_array[10340] <= 3'b101;
      memory_array[10341] <= 3'b101;
      memory_array[10342] <= 3'b111;
      memory_array[10343] <= 3'b110;
      memory_array[10344] <= 3'b110;
      memory_array[10345] <= 3'b000;
      memory_array[10346] <= 3'b000;
      memory_array[10347] <= 3'b000;
      memory_array[10348] <= 3'b110;
      memory_array[10349] <= 3'b110;
      memory_array[10350] <= 3'b101;
      memory_array[10351] <= 3'b101;
      memory_array[10352] <= 3'b101;
      memory_array[10353] <= 3'b101;
      memory_array[10354] <= 3'b101;
      memory_array[10355] <= 3'b101;
      memory_array[10356] <= 3'b101;
      memory_array[10357] <= 3'b101;
      memory_array[10358] <= 3'b101;
      memory_array[10359] <= 3'b101;
      memory_array[10360] <= 3'b101;
      memory_array[10361] <= 3'b000;
      memory_array[10362] <= 3'b111;
      memory_array[10363] <= 3'b111;
      memory_array[10364] <= 3'b111;
      memory_array[10365] <= 3'b111;
      memory_array[10366] <= 3'b000;
      memory_array[10367] <= 3'b000;
      memory_array[10368] <= 3'b000;
      memory_array[10369] <= 3'b110;
      memory_array[10370] <= 3'b000;
      memory_array[10371] <= 3'b000;
      memory_array[10372] <= 3'b101;
      memory_array[10373] <= 3'b101;
      memory_array[10374] <= 3'b000;
      memory_array[10375] <= 3'b000;
      memory_array[10376] <= 3'b000;
      memory_array[10377] <= 3'b000;
      memory_array[10378] <= 3'b110;
      memory_array[10379] <= 3'b110;
      memory_array[10380] <= 3'b000;
      memory_array[10381] <= 3'b000;
      memory_array[10382] <= 3'b000;
      memory_array[10383] <= 3'b110;
      memory_array[10384] <= 3'b110;
      memory_array[10385] <= 3'b000;
      memory_array[10386] <= 3'b101;
      memory_array[10387] <= 3'b000;
      memory_array[10388] <= 3'b110;
      memory_array[10389] <= 3'b000;
      memory_array[10390] <= 3'b000;
      memory_array[10391] <= 3'b101;
      memory_array[10392] <= 3'b101;
      memory_array[10393] <= 3'b101;
      memory_array[10394] <= 3'b101;
      memory_array[10395] <= 3'b111;
      memory_array[10396] <= 3'b111;
      memory_array[10397] <= 3'b101;
      memory_array[10398] <= 3'b101;
      memory_array[10399] <= 3'b101;
      memory_array[10400] <= 3'b101;
      memory_array[10401] <= 3'b101;
      memory_array[10402] <= 3'b101;
      memory_array[10403] <= 3'b101;
      memory_array[10404] <= 3'b101;
      memory_array[10405] <= 3'b101;
      memory_array[10406] <= 3'b101;
      memory_array[10407] <= 3'b101;
      memory_array[10408] <= 3'b101;
      memory_array[10409] <= 3'b000;
      memory_array[10410] <= 3'b000;
      memory_array[10411] <= 3'b000;
      memory_array[10412] <= 3'b000;
      memory_array[10413] <= 3'b101;
      memory_array[10414] <= 3'b101;
      memory_array[10415] <= 3'b000;
      memory_array[10416] <= 3'b000;
      memory_array[10417] <= 3'b000;
      memory_array[10418] <= 3'b110;
      memory_array[10419] <= 3'b000;
      memory_array[10420] <= 3'b000;
      memory_array[10421] <= 3'b000;
      memory_array[10422] <= 3'b000;
      memory_array[10423] <= 3'b110;
      memory_array[10424] <= 3'b111;
      memory_array[10425] <= 3'b000;
      memory_array[10426] <= 3'b101;
      memory_array[10427] <= 3'b000;
      memory_array[10428] <= 3'b101;
      memory_array[10429] <= 3'b110;
      memory_array[10430] <= 3'b000;
      memory_array[10431] <= 3'b000;
      memory_array[10432] <= 3'b000;
      memory_array[10433] <= 3'b000;
      memory_array[10434] <= 3'b111;
      memory_array[10435] <= 3'b111;
      memory_array[10436] <= 3'b111;
      memory_array[10437] <= 3'b111;
      memory_array[10438] <= 3'b000;
      memory_array[10439] <= 3'b101;
      memory_array[10440] <= 3'b101;
      memory_array[10441] <= 3'b101;
      memory_array[10442] <= 3'b101;
      memory_array[10443] <= 3'b101;
      memory_array[10444] <= 3'b101;
      memory_array[10445] <= 3'b101;
      memory_array[10446] <= 3'b101;
      memory_array[10447] <= 3'b101;
      memory_array[10448] <= 3'b101;
      memory_array[10449] <= 3'b101;
      memory_array[10450] <= 3'b101;
      memory_array[10451] <= 3'b101;
      memory_array[10452] <= 3'b101;
      memory_array[10453] <= 3'b101;
      memory_array[10454] <= 3'b101;
      memory_array[10455] <= 3'b101;
      memory_array[10456] <= 3'b101;
      memory_array[10457] <= 3'b101;
      memory_array[10458] <= 3'b101;
      memory_array[10459] <= 3'b101;
      memory_array[10460] <= 3'b101;
      memory_array[10461] <= 3'b101;
      memory_array[10462] <= 3'b101;
      memory_array[10463] <= 3'b101;
      memory_array[10464] <= 3'b101;
      memory_array[10465] <= 3'b101;
      memory_array[10466] <= 3'b101;
      memory_array[10467] <= 3'b000;
      memory_array[10468] <= 3'b101;
      memory_array[10469] <= 3'b101;
      memory_array[10470] <= 3'b101;
      memory_array[10471] <= 3'b101;
      memory_array[10472] <= 3'b000;
      memory_array[10473] <= 3'b111;
      memory_array[10474] <= 3'b101;
      memory_array[10475] <= 3'b000;
      memory_array[10476] <= 3'b000;
      memory_array[10477] <= 3'b101;
      memory_array[10478] <= 3'b101;
      memory_array[10479] <= 3'b101;
      memory_array[10480] <= 3'b000;
      memory_array[10481] <= 3'b111;
      memory_array[10482] <= 3'b101;
      memory_array[10483] <= 3'b111;
      memory_array[10484] <= 3'b111;
      memory_array[10485] <= 3'b111;
      memory_array[10486] <= 3'b101;
      memory_array[10487] <= 3'b101;
      memory_array[10488] <= 3'b111;
      memory_array[10489] <= 3'b111;
      memory_array[10490] <= 3'b111;
      memory_array[10491] <= 3'b101;
      memory_array[10492] <= 3'b000;
      memory_array[10493] <= 3'b111;
      memory_array[10494] <= 3'b111;
      memory_array[10495] <= 3'b111;
      memory_array[10496] <= 3'b111;
      memory_array[10497] <= 3'b111;
      memory_array[10498] <= 3'b111;
      memory_array[10499] <= 3'b111;
      memory_array[10500] <= 3'b111;
      memory_array[10501] <= 3'b111;
      memory_array[10502] <= 3'b111;
      memory_array[10503] <= 3'b111;
      memory_array[10504] <= 3'b101;
      memory_array[10505] <= 3'b111;
      memory_array[10506] <= 3'b000;
      memory_array[10507] <= 3'b110;
      memory_array[10508] <= 3'b110;
      memory_array[10509] <= 3'b110;
      memory_array[10510] <= 3'b000;
      memory_array[10511] <= 3'b101;
      memory_array[10512] <= 3'b101;
      memory_array[10513] <= 3'b101;
      memory_array[10514] <= 3'b101;
      memory_array[10515] <= 3'b101;
      memory_array[10516] <= 3'b101;
      memory_array[10517] <= 3'b101;
      memory_array[10518] <= 3'b111;
      memory_array[10519] <= 3'b000;
      memory_array[10520] <= 3'b101;
      memory_array[10521] <= 3'b101;
      memory_array[10522] <= 3'b101;
      memory_array[10523] <= 3'b101;
      memory_array[10524] <= 3'b101;
      memory_array[10525] <= 3'b101;
      memory_array[10526] <= 3'b101;
      memory_array[10527] <= 3'b101;
      memory_array[10528] <= 3'b101;
      memory_array[10529] <= 3'b110;
      memory_array[10530] <= 3'b110;
      memory_array[10531] <= 3'b110;
      memory_array[10532] <= 3'b000;
      memory_array[10533] <= 3'b110;
      memory_array[10534] <= 3'b110;
      memory_array[10535] <= 3'b110;
      memory_array[10536] <= 3'b101;
      memory_array[10537] <= 3'b101;
      memory_array[10538] <= 3'b110;
      memory_array[10539] <= 3'b110;
      memory_array[10540] <= 3'b110;
      memory_array[10541] <= 3'b000;
      memory_array[10542] <= 3'b101;
      memory_array[10543] <= 3'b101;
      memory_array[10544] <= 3'b110;
      memory_array[10545] <= 3'b111;
      memory_array[10546] <= 3'b101;
      memory_array[10547] <= 3'b101;
      memory_array[10548] <= 3'b110;
      memory_array[10549] <= 3'b101;
      memory_array[10550] <= 3'b101;
      memory_array[10551] <= 3'b101;
      memory_array[10552] <= 3'b101;
      memory_array[10553] <= 3'b101;
      memory_array[10554] <= 3'b101;
      memory_array[10555] <= 3'b101;
      memory_array[10556] <= 3'b101;
      memory_array[10557] <= 3'b101;
      memory_array[10558] <= 3'b101;
      memory_array[10559] <= 3'b101;
      memory_array[10560] <= 3'b101;
      memory_array[10561] <= 3'b000;
      memory_array[10562] <= 3'b111;
      memory_array[10563] <= 3'b111;
      memory_array[10564] <= 3'b111;
      memory_array[10565] <= 3'b111;
      memory_array[10566] <= 3'b000;
      memory_array[10567] <= 3'b000;
      memory_array[10568] <= 3'b110;
      memory_array[10569] <= 3'b110;
      memory_array[10570] <= 3'b000;
      memory_array[10571] <= 3'b101;
      memory_array[10572] <= 3'b000;
      memory_array[10573] <= 3'b101;
      memory_array[10574] <= 3'b101;
      memory_array[10575] <= 3'b111;
      memory_array[10576] <= 3'b000;
      memory_array[10577] <= 3'b000;
      memory_array[10578] <= 3'b110;
      memory_array[10579] <= 3'b000;
      memory_array[10580] <= 3'b000;
      memory_array[10581] <= 3'b000;
      memory_array[10582] <= 3'b101;
      memory_array[10583] <= 3'b000;
      memory_array[10584] <= 3'b000;
      memory_array[10585] <= 3'b101;
      memory_array[10586] <= 3'b101;
      memory_array[10587] <= 3'b000;
      memory_array[10588] <= 3'b110;
      memory_array[10589] <= 3'b000;
      memory_array[10590] <= 3'b000;
      memory_array[10591] <= 3'b101;
      memory_array[10592] <= 3'b111;
      memory_array[10593] <= 3'b101;
      memory_array[10594] <= 3'b101;
      memory_array[10595] <= 3'b101;
      memory_array[10596] <= 3'b101;
      memory_array[10597] <= 3'b101;
      memory_array[10598] <= 3'b101;
      memory_array[10599] <= 3'b101;
      memory_array[10600] <= 3'b101;
      memory_array[10601] <= 3'b101;
      memory_array[10602] <= 3'b101;
      memory_array[10603] <= 3'b101;
      memory_array[10604] <= 3'b101;
      memory_array[10605] <= 3'b101;
      memory_array[10606] <= 3'b101;
      memory_array[10607] <= 3'b101;
      memory_array[10608] <= 3'b101;
      memory_array[10609] <= 3'b000;
      memory_array[10610] <= 3'b000;
      memory_array[10611] <= 3'b101;
      memory_array[10612] <= 3'b000;
      memory_array[10613] <= 3'b000;
      memory_array[10614] <= 3'b000;
      memory_array[10615] <= 3'b000;
      memory_array[10616] <= 3'b000;
      memory_array[10617] <= 3'b101;
      memory_array[10618] <= 3'b000;
      memory_array[10619] <= 3'b000;
      memory_array[10620] <= 3'b110;
      memory_array[10621] <= 3'b110;
      memory_array[10622] <= 3'b110;
      memory_array[10623] <= 3'b000;
      memory_array[10624] <= 3'b111;
      memory_array[10625] <= 3'b110;
      memory_array[10626] <= 3'b000;
      memory_array[10627] <= 3'b101;
      memory_array[10628] <= 3'b101;
      memory_array[10629] <= 3'b000;
      memory_array[10630] <= 3'b110;
      memory_array[10631] <= 3'b110;
      memory_array[10632] <= 3'b110;
      memory_array[10633] <= 3'b000;
      memory_array[10634] <= 3'b111;
      memory_array[10635] <= 3'b111;
      memory_array[10636] <= 3'b111;
      memory_array[10637] <= 3'b111;
      memory_array[10638] <= 3'b000;
      memory_array[10639] <= 3'b101;
      memory_array[10640] <= 3'b101;
      memory_array[10641] <= 3'b101;
      memory_array[10642] <= 3'b101;
      memory_array[10643] <= 3'b101;
      memory_array[10644] <= 3'b101;
      memory_array[10645] <= 3'b101;
      memory_array[10646] <= 3'b101;
      memory_array[10647] <= 3'b101;
      memory_array[10648] <= 3'b101;
      memory_array[10649] <= 3'b101;
      memory_array[10650] <= 3'b101;
      memory_array[10651] <= 3'b101;
      memory_array[10652] <= 3'b101;
      memory_array[10653] <= 3'b101;
      memory_array[10654] <= 3'b101;
      memory_array[10655] <= 3'b101;
      memory_array[10656] <= 3'b101;
      memory_array[10657] <= 3'b101;
      memory_array[10658] <= 3'b101;
      memory_array[10659] <= 3'b101;
      memory_array[10660] <= 3'b101;
      memory_array[10661] <= 3'b101;
      memory_array[10662] <= 3'b101;
      memory_array[10663] <= 3'b101;
      memory_array[10664] <= 3'b101;
      memory_array[10665] <= 3'b101;
      memory_array[10666] <= 3'b101;
      memory_array[10667] <= 3'b101;
      memory_array[10668] <= 3'b000;
      memory_array[10669] <= 3'b101;
      memory_array[10670] <= 3'b101;
      memory_array[10671] <= 3'b101;
      memory_array[10672] <= 3'b000;
      memory_array[10673] <= 3'b111;
      memory_array[10674] <= 3'b000;
      memory_array[10675] <= 3'b101;
      memory_array[10676] <= 3'b101;
      memory_array[10677] <= 3'b000;
      memory_array[10678] <= 3'b000;
      memory_array[10679] <= 3'b000;
      memory_array[10680] <= 3'b000;
      memory_array[10681] <= 3'b111;
      memory_array[10682] <= 3'b101;
      memory_array[10683] <= 3'b111;
      memory_array[10684] <= 3'b111;
      memory_array[10685] <= 3'b111;
      memory_array[10686] <= 3'b101;
      memory_array[10687] <= 3'b111;
      memory_array[10688] <= 3'b111;
      memory_array[10689] <= 3'b111;
      memory_array[10690] <= 3'b111;
      memory_array[10691] <= 3'b111;
      memory_array[10692] <= 3'b000;
      memory_array[10693] <= 3'b000;
      memory_array[10694] <= 3'b111;
      memory_array[10695] <= 3'b111;
      memory_array[10696] <= 3'b101;
      memory_array[10697] <= 3'b111;
      memory_array[10698] <= 3'b111;
      memory_array[10699] <= 3'b000;
      memory_array[10700] <= 3'b101;
      memory_array[10701] <= 3'b111;
      memory_array[10702] <= 3'b111;
      memory_array[10703] <= 3'b111;
      memory_array[10704] <= 3'b000;
      memory_array[10705] <= 3'b101;
      memory_array[10706] <= 3'b111;
      memory_array[10707] <= 3'b101;
      memory_array[10708] <= 3'b000;
      memory_array[10709] <= 3'b000;
      memory_array[10710] <= 3'b000;
      memory_array[10711] <= 3'b101;
      memory_array[10712] <= 3'b101;
      memory_array[10713] <= 3'b101;
      memory_array[10714] <= 3'b101;
      memory_array[10715] <= 3'b101;
      memory_array[10716] <= 3'b101;
      memory_array[10717] <= 3'b101;
      memory_array[10718] <= 3'b111;
      memory_array[10719] <= 3'b000;
      memory_array[10720] <= 3'b101;
      memory_array[10721] <= 3'b101;
      memory_array[10722] <= 3'b101;
      memory_array[10723] <= 3'b101;
      memory_array[10724] <= 3'b101;
      memory_array[10725] <= 3'b101;
      memory_array[10726] <= 3'b101;
      memory_array[10727] <= 3'b101;
      memory_array[10728] <= 3'b101;
      memory_array[10729] <= 3'b101;
      memory_array[10730] <= 3'b101;
      memory_array[10731] <= 3'b110;
      memory_array[10732] <= 3'b110;
      memory_array[10733] <= 3'b000;
      memory_array[10734] <= 3'b110;
      memory_array[10735] <= 3'b110;
      memory_array[10736] <= 3'b110;
      memory_array[10737] <= 3'b101;
      memory_array[10738] <= 3'b101;
      memory_array[10739] <= 3'b101;
      memory_array[10740] <= 3'b110;
      memory_array[10741] <= 3'b110;
      memory_array[10742] <= 3'b110;
      memory_array[10743] <= 3'b101;
      memory_array[10744] <= 3'b000;
      memory_array[10745] <= 3'b101;
      memory_array[10746] <= 3'b110;
      memory_array[10747] <= 3'b101;
      memory_array[10748] <= 3'b101;
      memory_array[10749] <= 3'b101;
      memory_array[10750] <= 3'b101;
      memory_array[10751] <= 3'b101;
      memory_array[10752] <= 3'b101;
      memory_array[10753] <= 3'b101;
      memory_array[10754] <= 3'b101;
      memory_array[10755] <= 3'b101;
      memory_array[10756] <= 3'b101;
      memory_array[10757] <= 3'b101;
      memory_array[10758] <= 3'b101;
      memory_array[10759] <= 3'b101;
      memory_array[10760] <= 3'b101;
      memory_array[10761] <= 3'b000;
      memory_array[10762] <= 3'b111;
      memory_array[10763] <= 3'b111;
      memory_array[10764] <= 3'b111;
      memory_array[10765] <= 3'b111;
      memory_array[10766] <= 3'b000;
      memory_array[10767] <= 3'b110;
      memory_array[10768] <= 3'b000;
      memory_array[10769] <= 3'b000;
      memory_array[10770] <= 3'b110;
      memory_array[10771] <= 3'b101;
      memory_array[10772] <= 3'b101;
      memory_array[10773] <= 3'b000;
      memory_array[10774] <= 3'b111;
      memory_array[10775] <= 3'b111;
      memory_array[10776] <= 3'b110;
      memory_array[10777] <= 3'b110;
      memory_array[10778] <= 3'b000;
      memory_array[10779] <= 3'b000;
      memory_array[10780] <= 3'b000;
      memory_array[10781] <= 3'b000;
      memory_array[10782] <= 3'b000;
      memory_array[10783] <= 3'b000;
      memory_array[10784] <= 3'b000;
      memory_array[10785] <= 3'b000;
      memory_array[10786] <= 3'b000;
      memory_array[10787] <= 3'b101;
      memory_array[10788] <= 3'b101;
      memory_array[10789] <= 3'b000;
      memory_array[10790] <= 3'b000;
      memory_array[10791] <= 3'b101;
      memory_array[10792] <= 3'b101;
      memory_array[10793] <= 3'b101;
      memory_array[10794] <= 3'b101;
      memory_array[10795] <= 3'b101;
      memory_array[10796] <= 3'b101;
      memory_array[10797] <= 3'b101;
      memory_array[10798] <= 3'b101;
      memory_array[10799] <= 3'b101;
      memory_array[10800] <= 3'b101;
      memory_array[10801] <= 3'b101;
      memory_array[10802] <= 3'b101;
      memory_array[10803] <= 3'b111;
      memory_array[10804] <= 3'b111;
      memory_array[10805] <= 3'b101;
      memory_array[10806] <= 3'b101;
      memory_array[10807] <= 3'b101;
      memory_array[10808] <= 3'b101;
      memory_array[10809] <= 3'b000;
      memory_array[10810] <= 3'b000;
      memory_array[10811] <= 3'b000;
      memory_array[10812] <= 3'b101;
      memory_array[10813] <= 3'b000;
      memory_array[10814] <= 3'b110;
      memory_array[10815] <= 3'b000;
      memory_array[10816] <= 3'b000;
      memory_array[10817] <= 3'b000;
      memory_array[10818] <= 3'b000;
      memory_array[10819] <= 3'b110;
      memory_array[10820] <= 3'b000;
      memory_array[10821] <= 3'b000;
      memory_array[10822] <= 3'b000;
      memory_array[10823] <= 3'b110;
      memory_array[10824] <= 3'b111;
      memory_array[10825] <= 3'b000;
      memory_array[10826] <= 3'b101;
      memory_array[10827] <= 3'b000;
      memory_array[10828] <= 3'b101;
      memory_array[10829] <= 3'b110;
      memory_array[10830] <= 3'b000;
      memory_array[10831] <= 3'b000;
      memory_array[10832] <= 3'b000;
      memory_array[10833] <= 3'b000;
      memory_array[10834] <= 3'b111;
      memory_array[10835] <= 3'b111;
      memory_array[10836] <= 3'b111;
      memory_array[10837] <= 3'b111;
      memory_array[10838] <= 3'b000;
      memory_array[10839] <= 3'b101;
      memory_array[10840] <= 3'b101;
      memory_array[10841] <= 3'b101;
      memory_array[10842] <= 3'b101;
      memory_array[10843] <= 3'b101;
      memory_array[10844] <= 3'b101;
      memory_array[10845] <= 3'b101;
      memory_array[10846] <= 3'b101;
      memory_array[10847] <= 3'b101;
      memory_array[10848] <= 3'b101;
      memory_array[10849] <= 3'b101;
      memory_array[10850] <= 3'b101;
      memory_array[10851] <= 3'b101;
      memory_array[10852] <= 3'b101;
      memory_array[10853] <= 3'b101;
      memory_array[10854] <= 3'b101;
      memory_array[10855] <= 3'b101;
      memory_array[10856] <= 3'b101;
      memory_array[10857] <= 3'b101;
      memory_array[10858] <= 3'b101;
      memory_array[10859] <= 3'b101;
      memory_array[10860] <= 3'b101;
      memory_array[10861] <= 3'b101;
      memory_array[10862] <= 3'b101;
      memory_array[10863] <= 3'b101;
      memory_array[10864] <= 3'b101;
      memory_array[10865] <= 3'b101;
      memory_array[10866] <= 3'b000;
      memory_array[10867] <= 3'b111;
      memory_array[10868] <= 3'b101;
      memory_array[10869] <= 3'b101;
      memory_array[10870] <= 3'b101;
      memory_array[10871] <= 3'b101;
      memory_array[10872] <= 3'b000;
      memory_array[10873] <= 3'b101;
      memory_array[10874] <= 3'b111;
      memory_array[10875] <= 3'b111;
      memory_array[10876] <= 3'b111;
      memory_array[10877] <= 3'b111;
      memory_array[10878] <= 3'b101;
      memory_array[10879] <= 3'b101;
      memory_array[10880] <= 3'b000;
      memory_array[10881] <= 3'b111;
      memory_array[10882] <= 3'b101;
      memory_array[10883] <= 3'b111;
      memory_array[10884] <= 3'b111;
      memory_array[10885] <= 3'b111;
      memory_array[10886] <= 3'b101;
      memory_array[10887] <= 3'b111;
      memory_array[10888] <= 3'b111;
      memory_array[10889] <= 3'b111;
      memory_array[10890] <= 3'b111;
      memory_array[10891] <= 3'b111;
      memory_array[10892] <= 3'b000;
      memory_array[10893] <= 3'b101;
      memory_array[10894] <= 3'b111;
      memory_array[10895] <= 3'b111;
      memory_array[10896] <= 3'b000;
      memory_array[10897] <= 3'b111;
      memory_array[10898] <= 3'b111;
      memory_array[10899] <= 3'b101;
      memory_array[10900] <= 3'b000;
      memory_array[10901] <= 3'b111;
      memory_array[10902] <= 3'b111;
      memory_array[10903] <= 3'b111;
      memory_array[10904] <= 3'b000;
      memory_array[10905] <= 3'b000;
      memory_array[10906] <= 3'b111;
      memory_array[10907] <= 3'b000;
      memory_array[10908] <= 3'b000;
      memory_array[10909] <= 3'b101;
      memory_array[10910] <= 3'b000;
      memory_array[10911] <= 3'b101;
      memory_array[10912] <= 3'b101;
      memory_array[10913] <= 3'b101;
      memory_array[10914] <= 3'b101;
      memory_array[10915] <= 3'b101;
      memory_array[10916] <= 3'b101;
      memory_array[10917] <= 3'b101;
      memory_array[10918] <= 3'b111;
      memory_array[10919] <= 3'b000;
      memory_array[10920] <= 3'b101;
      memory_array[10921] <= 3'b101;
      memory_array[10922] <= 3'b101;
      memory_array[10923] <= 3'b101;
      memory_array[10924] <= 3'b101;
      memory_array[10925] <= 3'b101;
      memory_array[10926] <= 3'b101;
      memory_array[10927] <= 3'b101;
      memory_array[10928] <= 3'b101;
      memory_array[10929] <= 3'b101;
      memory_array[10930] <= 3'b101;
      memory_array[10931] <= 3'b101;
      memory_array[10932] <= 3'b101;
      memory_array[10933] <= 3'b110;
      memory_array[10934] <= 3'b101;
      memory_array[10935] <= 3'b000;
      memory_array[10936] <= 3'b101;
      memory_array[10937] <= 3'b101;
      memory_array[10938] <= 3'b101;
      memory_array[10939] <= 3'b110;
      memory_array[10940] <= 3'b101;
      memory_array[10941] <= 3'b000;
      memory_array[10942] <= 3'b101;
      memory_array[10943] <= 3'b101;
      memory_array[10944] <= 3'b110;
      memory_array[10945] <= 3'b101;
      memory_array[10946] <= 3'b101;
      memory_array[10947] <= 3'b101;
      memory_array[10948] <= 3'b101;
      memory_array[10949] <= 3'b101;
      memory_array[10950] <= 3'b101;
      memory_array[10951] <= 3'b101;
      memory_array[10952] <= 3'b101;
      memory_array[10953] <= 3'b101;
      memory_array[10954] <= 3'b101;
      memory_array[10955] <= 3'b101;
      memory_array[10956] <= 3'b101;
      memory_array[10957] <= 3'b101;
      memory_array[10958] <= 3'b101;
      memory_array[10959] <= 3'b101;
      memory_array[10960] <= 3'b101;
      memory_array[10961] <= 3'b000;
      memory_array[10962] <= 3'b111;
      memory_array[10963] <= 3'b111;
      memory_array[10964] <= 3'b111;
      memory_array[10965] <= 3'b111;
      memory_array[10966] <= 3'b000;
      memory_array[10967] <= 3'b000;
      memory_array[10968] <= 3'b110;
      memory_array[10969] <= 3'b110;
      memory_array[10970] <= 3'b000;
      memory_array[10971] <= 3'b101;
      memory_array[10972] <= 3'b000;
      memory_array[10973] <= 3'b101;
      memory_array[10974] <= 3'b101;
      memory_array[10975] <= 3'b111;
      memory_array[10976] <= 3'b000;
      memory_array[10977] <= 3'b000;
      memory_array[10978] <= 3'b110;
      memory_array[10979] <= 3'b110;
      memory_array[10980] <= 3'b000;
      memory_array[10981] <= 3'b000;
      memory_array[10982] <= 3'b000;
      memory_array[10983] <= 3'b110;
      memory_array[10984] <= 3'b110;
      memory_array[10985] <= 3'b000;
      memory_array[10986] <= 3'b000;
      memory_array[10987] <= 3'b000;
      memory_array[10988] <= 3'b000;
      memory_array[10989] <= 3'b000;
      memory_array[10990] <= 3'b000;
      memory_array[10991] <= 3'b101;
      memory_array[10992] <= 3'b101;
      memory_array[10993] <= 3'b101;
      memory_array[10994] <= 3'b101;
      memory_array[10995] <= 3'b111;
      memory_array[10996] <= 3'b111;
      memory_array[10997] <= 3'b101;
      memory_array[10998] <= 3'b101;
      memory_array[10999] <= 3'b101;
      memory_array[11000] <= 3'b101;
      memory_array[11001] <= 3'b101;
      memory_array[11002] <= 3'b110;
      memory_array[11003] <= 3'b101;
      memory_array[11004] <= 3'b101;
      memory_array[11005] <= 3'b110;
      memory_array[11006] <= 3'b101;
      memory_array[11007] <= 3'b101;
      memory_array[11008] <= 3'b101;
      memory_array[11009] <= 3'b000;
      memory_array[11010] <= 3'b000;
      memory_array[11011] <= 3'b110;
      memory_array[11012] <= 3'b000;
      memory_array[11013] <= 3'b101;
      memory_array[11014] <= 3'b000;
      memory_array[11015] <= 3'b110;
      memory_array[11016] <= 3'b110;
      memory_array[11017] <= 3'b110;
      memory_array[11018] <= 3'b000;
      memory_array[11019] <= 3'b000;
      memory_array[11020] <= 3'b110;
      memory_array[11021] <= 3'b110;
      memory_array[11022] <= 3'b110;
      memory_array[11023] <= 3'b000;
      memory_array[11024] <= 3'b000;
      memory_array[11025] <= 3'b110;
      memory_array[11026] <= 3'b101;
      memory_array[11027] <= 3'b000;
      memory_array[11028] <= 3'b000;
      memory_array[11029] <= 3'b000;
      memory_array[11030] <= 3'b110;
      memory_array[11031] <= 3'b110;
      memory_array[11032] <= 3'b110;
      memory_array[11033] <= 3'b000;
      memory_array[11034] <= 3'b111;
      memory_array[11035] <= 3'b111;
      memory_array[11036] <= 3'b111;
      memory_array[11037] <= 3'b111;
      memory_array[11038] <= 3'b000;
      memory_array[11039] <= 3'b101;
      memory_array[11040] <= 3'b101;
      memory_array[11041] <= 3'b101;
      memory_array[11042] <= 3'b101;
      memory_array[11043] <= 3'b101;
      memory_array[11044] <= 3'b101;
      memory_array[11045] <= 3'b101;
      memory_array[11046] <= 3'b101;
      memory_array[11047] <= 3'b101;
      memory_array[11048] <= 3'b101;
      memory_array[11049] <= 3'b101;
      memory_array[11050] <= 3'b101;
      memory_array[11051] <= 3'b101;
      memory_array[11052] <= 3'b101;
      memory_array[11053] <= 3'b101;
      memory_array[11054] <= 3'b101;
      memory_array[11055] <= 3'b101;
      memory_array[11056] <= 3'b101;
      memory_array[11057] <= 3'b101;
      memory_array[11058] <= 3'b101;
      memory_array[11059] <= 3'b101;
      memory_array[11060] <= 3'b101;
      memory_array[11061] <= 3'b101;
      memory_array[11062] <= 3'b101;
      memory_array[11063] <= 3'b101;
      memory_array[11064] <= 3'b101;
      memory_array[11065] <= 3'b101;
      memory_array[11066] <= 3'b101;
      memory_array[11067] <= 3'b111;
      memory_array[11068] <= 3'b111;
      memory_array[11069] <= 3'b101;
      memory_array[11070] <= 3'b101;
      memory_array[11071] <= 3'b101;
      memory_array[11072] <= 3'b000;
      memory_array[11073] <= 3'b000;
      memory_array[11074] <= 3'b111;
      memory_array[11075] <= 3'b111;
      memory_array[11076] <= 3'b101;
      memory_array[11077] <= 3'b111;
      memory_array[11078] <= 3'b101;
      memory_array[11079] <= 3'b101;
      memory_array[11080] <= 3'b101;
      memory_array[11081] <= 3'b101;
      memory_array[11082] <= 3'b101;
      memory_array[11083] <= 3'b101;
      memory_array[11084] <= 3'b101;
      memory_array[11085] <= 3'b000;
      memory_array[11086] <= 3'b000;
      memory_array[11087] <= 3'b101;
      memory_array[11088] <= 3'b111;
      memory_array[11089] <= 3'b111;
      memory_array[11090] <= 3'b111;
      memory_array[11091] <= 3'b111;
      memory_array[11092] <= 3'b000;
      memory_array[11093] <= 3'b000;
      memory_array[11094] <= 3'b111;
      memory_array[11095] <= 3'b111;
      memory_array[11096] <= 3'b101;
      memory_array[11097] <= 3'b111;
      memory_array[11098] <= 3'b111;
      memory_array[11099] <= 3'b000;
      memory_array[11100] <= 3'b101;
      memory_array[11101] <= 3'b111;
      memory_array[11102] <= 3'b111;
      memory_array[11103] <= 3'b111;
      memory_array[11104] <= 3'b000;
      memory_array[11105] <= 3'b101;
      memory_array[11106] <= 3'b111;
      memory_array[11107] <= 3'b101;
      memory_array[11108] <= 3'b000;
      memory_array[11109] <= 3'b000;
      memory_array[11110] <= 3'b101;
      memory_array[11111] <= 3'b000;
      memory_array[11112] <= 3'b101;
      memory_array[11113] <= 3'b101;
      memory_array[11114] <= 3'b101;
      memory_array[11115] <= 3'b101;
      memory_array[11116] <= 3'b101;
      memory_array[11117] <= 3'b101;
      memory_array[11118] <= 3'b111;
      memory_array[11119] <= 3'b000;
      memory_array[11120] <= 3'b101;
      memory_array[11121] <= 3'b101;
      memory_array[11122] <= 3'b101;
      memory_array[11123] <= 3'b101;
      memory_array[11124] <= 3'b101;
      memory_array[11125] <= 3'b101;
      memory_array[11126] <= 3'b101;
      memory_array[11127] <= 3'b101;
      memory_array[11128] <= 3'b101;
      memory_array[11129] <= 3'b101;
      memory_array[11130] <= 3'b101;
      memory_array[11131] <= 3'b101;
      memory_array[11132] <= 3'b101;
      memory_array[11133] <= 3'b000;
      memory_array[11134] <= 3'b101;
      memory_array[11135] <= 3'b101;
      memory_array[11136] <= 3'b101;
      memory_array[11137] <= 3'b101;
      memory_array[11138] <= 3'b101;
      memory_array[11139] <= 3'b101;
      memory_array[11140] <= 3'b101;
      memory_array[11141] <= 3'b110;
      memory_array[11142] <= 3'b101;
      memory_array[11143] <= 3'b101;
      memory_array[11144] <= 3'b110;
      memory_array[11145] <= 3'b101;
      memory_array[11146] <= 3'b101;
      memory_array[11147] <= 3'b101;
      memory_array[11148] <= 3'b101;
      memory_array[11149] <= 3'b101;
      memory_array[11150] <= 3'b101;
      memory_array[11151] <= 3'b101;
      memory_array[11152] <= 3'b101;
      memory_array[11153] <= 3'b101;
      memory_array[11154] <= 3'b101;
      memory_array[11155] <= 3'b101;
      memory_array[11156] <= 3'b101;
      memory_array[11157] <= 3'b101;
      memory_array[11158] <= 3'b101;
      memory_array[11159] <= 3'b101;
      memory_array[11160] <= 3'b101;
      memory_array[11161] <= 3'b000;
      memory_array[11162] <= 3'b111;
      memory_array[11163] <= 3'b111;
      memory_array[11164] <= 3'b111;
      memory_array[11165] <= 3'b111;
      memory_array[11166] <= 3'b000;
      memory_array[11167] <= 3'b110;
      memory_array[11168] <= 3'b000;
      memory_array[11169] <= 3'b000;
      memory_array[11170] <= 3'b110;
      memory_array[11171] <= 3'b110;
      memory_array[11172] <= 3'b000;
      memory_array[11173] <= 3'b101;
      memory_array[11174] <= 3'b000;
      memory_array[11175] <= 3'b000;
      memory_array[11176] <= 3'b110;
      memory_array[11177] <= 3'b110;
      memory_array[11178] <= 3'b000;
      memory_array[11179] <= 3'b000;
      memory_array[11180] <= 3'b110;
      memory_array[11181] <= 3'b110;
      memory_array[11182] <= 3'b110;
      memory_array[11183] <= 3'b000;
      memory_array[11184] <= 3'b000;
      memory_array[11185] <= 3'b110;
      memory_array[11186] <= 3'b101;
      memory_array[11187] <= 3'b000;
      memory_array[11188] <= 3'b000;
      memory_array[11189] <= 3'b000;
      memory_array[11190] <= 3'b000;
      memory_array[11191] <= 3'b101;
      memory_array[11192] <= 3'b101;
      memory_array[11193] <= 3'b101;
      memory_array[11194] <= 3'b000;
      memory_array[11195] <= 3'b101;
      memory_array[11196] <= 3'b101;
      memory_array[11197] <= 3'b110;
      memory_array[11198] <= 3'b101;
      memory_array[11199] <= 3'b101;
      memory_array[11200] <= 3'b101;
      memory_array[11201] <= 3'b110;
      memory_array[11202] <= 3'b110;
      memory_array[11203] <= 3'b000;
      memory_array[11204] <= 3'b000;
      memory_array[11205] <= 3'b110;
      memory_array[11206] <= 3'b110;
      memory_array[11207] <= 3'b101;
      memory_array[11208] <= 3'b101;
      memory_array[11209] <= 3'b000;
      memory_array[11210] <= 3'b000;
      memory_array[11211] <= 3'b110;
      memory_array[11212] <= 3'b000;
      memory_array[11213] <= 3'b000;
      memory_array[11214] <= 3'b000;
      memory_array[11215] <= 3'b110;
      memory_array[11216] <= 3'b110;
      memory_array[11217] <= 3'b110;
      memory_array[11218] <= 3'b000;
      memory_array[11219] <= 3'b000;
      memory_array[11220] <= 3'b000;
      memory_array[11221] <= 3'b101;
      memory_array[11222] <= 3'b101;
      memory_array[11223] <= 3'b000;
      memory_array[11224] <= 3'b000;
      memory_array[11225] <= 3'b000;
      memory_array[11226] <= 3'b000;
      memory_array[11227] <= 3'b110;
      memory_array[11228] <= 3'b000;
      memory_array[11229] <= 3'b000;
      memory_array[11230] <= 3'b101;
      memory_array[11231] <= 3'b101;
      memory_array[11232] <= 3'b101;
      memory_array[11233] <= 3'b000;
      memory_array[11234] <= 3'b111;
      memory_array[11235] <= 3'b111;
      memory_array[11236] <= 3'b111;
      memory_array[11237] <= 3'b111;
      memory_array[11238] <= 3'b101;
      memory_array[11239] <= 3'b101;
      memory_array[11240] <= 3'b101;
      memory_array[11241] <= 3'b101;
      memory_array[11242] <= 3'b101;
      memory_array[11243] <= 3'b101;
      memory_array[11244] <= 3'b101;
      memory_array[11245] <= 3'b101;
      memory_array[11246] <= 3'b101;
      memory_array[11247] <= 3'b101;
      memory_array[11248] <= 3'b101;
      memory_array[11249] <= 3'b101;
      memory_array[11250] <= 3'b101;
      memory_array[11251] <= 3'b101;
      memory_array[11252] <= 3'b101;
      memory_array[11253] <= 3'b101;
      memory_array[11254] <= 3'b000;
      memory_array[11255] <= 3'b000;
      memory_array[11256] <= 3'b000;
      memory_array[11257] <= 3'b101;
      memory_array[11258] <= 3'b000;
      memory_array[11259] <= 3'b101;
      memory_array[11260] <= 3'b101;
      memory_array[11261] <= 3'b101;
      memory_array[11262] <= 3'b101;
      memory_array[11263] <= 3'b101;
      memory_array[11264] <= 3'b101;
      memory_array[11265] <= 3'b101;
      memory_array[11266] <= 3'b111;
      memory_array[11267] <= 3'b111;
      memory_array[11268] <= 3'b111;
      memory_array[11269] <= 3'b101;
      memory_array[11270] <= 3'b101;
      memory_array[11271] <= 3'b101;
      memory_array[11272] <= 3'b111;
      memory_array[11273] <= 3'b101;
      memory_array[11274] <= 3'b101;
      memory_array[11275] <= 3'b101;
      memory_array[11276] <= 3'b101;
      memory_array[11277] <= 3'b101;
      memory_array[11278] <= 3'b000;
      memory_array[11279] <= 3'b000;
      memory_array[11280] <= 3'b101;
      memory_array[11281] <= 3'b111;
      memory_array[11282] <= 3'b111;
      memory_array[11283] <= 3'b000;
      memory_array[11284] <= 3'b111;
      memory_array[11285] <= 3'b111;
      memory_array[11286] <= 3'b101;
      memory_array[11287] <= 3'b101;
      memory_array[11288] <= 3'b101;
      memory_array[11289] <= 3'b111;
      memory_array[11290] <= 3'b111;
      memory_array[11291] <= 3'b111;
      memory_array[11292] <= 3'b101;
      memory_array[11293] <= 3'b101;
      memory_array[11294] <= 3'b110;
      memory_array[11295] <= 3'b111;
      memory_array[11296] <= 3'b111;
      memory_array[11297] <= 3'b111;
      memory_array[11298] <= 3'b111;
      memory_array[11299] <= 3'b111;
      memory_array[11300] <= 3'b111;
      memory_array[11301] <= 3'b111;
      memory_array[11302] <= 3'b111;
      memory_array[11303] <= 3'b111;
      memory_array[11304] <= 3'b101;
      memory_array[11305] <= 3'b101;
      memory_array[11306] <= 3'b111;
      memory_array[11307] <= 3'b101;
      memory_array[11308] <= 3'b101;
      memory_array[11309] <= 3'b000;
      memory_array[11310] <= 3'b101;
      memory_array[11311] <= 3'b000;
      memory_array[11312] <= 3'b000;
      memory_array[11313] <= 3'b000;
      memory_array[11314] <= 3'b101;
      memory_array[11315] <= 3'b101;
      memory_array[11316] <= 3'b101;
      memory_array[11317] <= 3'b101;
      memory_array[11318] <= 3'b111;
      memory_array[11319] <= 3'b110;
      memory_array[11320] <= 3'b101;
      memory_array[11321] <= 3'b101;
      memory_array[11322] <= 3'b101;
      memory_array[11323] <= 3'b101;
      memory_array[11324] <= 3'b101;
      memory_array[11325] <= 3'b101;
      memory_array[11326] <= 3'b101;
      memory_array[11327] <= 3'b101;
      memory_array[11328] <= 3'b101;
      memory_array[11329] <= 3'b101;
      memory_array[11330] <= 3'b101;
      memory_array[11331] <= 3'b101;
      memory_array[11332] <= 3'b101;
      memory_array[11333] <= 3'b111;
      memory_array[11334] <= 3'b101;
      memory_array[11335] <= 3'b101;
      memory_array[11336] <= 3'b101;
      memory_array[11337] <= 3'b101;
      memory_array[11338] <= 3'b101;
      memory_array[11339] <= 3'b101;
      memory_array[11340] <= 3'b101;
      memory_array[11341] <= 3'b101;
      memory_array[11342] <= 3'b101;
      memory_array[11343] <= 3'b101;
      memory_array[11344] <= 3'b110;
      memory_array[11345] <= 3'b110;
      memory_array[11346] <= 3'b110;
      memory_array[11347] <= 3'b110;
      memory_array[11348] <= 3'b101;
      memory_array[11349] <= 3'b101;
      memory_array[11350] <= 3'b101;
      memory_array[11351] <= 3'b101;
      memory_array[11352] <= 3'b101;
      memory_array[11353] <= 3'b101;
      memory_array[11354] <= 3'b101;
      memory_array[11355] <= 3'b101;
      memory_array[11356] <= 3'b101;
      memory_array[11357] <= 3'b101;
      memory_array[11358] <= 3'b101;
      memory_array[11359] <= 3'b101;
      memory_array[11360] <= 3'b101;
      memory_array[11361] <= 3'b101;
      memory_array[11362] <= 3'b111;
      memory_array[11363] <= 3'b111;
      memory_array[11364] <= 3'b111;
      memory_array[11365] <= 3'b111;
      memory_array[11366] <= 3'b000;
      memory_array[11367] <= 3'b101;
      memory_array[11368] <= 3'b101;
      memory_array[11369] <= 3'b101;
      memory_array[11370] <= 3'b101;
      memory_array[11371] <= 3'b110;
      memory_array[11372] <= 3'b110;
      memory_array[11373] <= 3'b000;
      memory_array[11374] <= 3'b000;
      memory_array[11375] <= 3'b110;
      memory_array[11376] <= 3'b000;
      memory_array[11377] <= 3'b101;
      memory_array[11378] <= 3'b101;
      memory_array[11379] <= 3'b000;
      memory_array[11380] <= 3'b000;
      memory_array[11381] <= 3'b110;
      memory_array[11382] <= 3'b110;
      memory_array[11383] <= 3'b000;
      memory_array[11384] <= 3'b000;
      memory_array[11385] <= 3'b000;
      memory_array[11386] <= 3'b000;
      memory_array[11387] <= 3'b110;
      memory_array[11388] <= 3'b000;
      memory_array[11389] <= 3'b000;
      memory_array[11390] <= 3'b000;
      memory_array[11391] <= 3'b101;
      memory_array[11392] <= 3'b110;
      memory_array[11393] <= 3'b000;
      memory_array[11394] <= 3'b000;
      memory_array[11395] <= 3'b110;
      memory_array[11396] <= 3'b110;
      memory_array[11397] <= 3'b110;
      memory_array[11398] <= 3'b000;
      memory_array[11399] <= 3'b101;
      memory_array[11400] <= 3'b000;
      memory_array[11401] <= 3'b000;
      memory_array[11402] <= 3'b000;
      memory_array[11403] <= 3'b110;
      memory_array[11404] <= 3'b110;
      memory_array[11405] <= 3'b000;
      memory_array[11406] <= 3'b000;
      memory_array[11407] <= 3'b000;
      memory_array[11408] <= 3'b101;
      memory_array[11409] <= 3'b000;
      memory_array[11410] <= 3'b000;
      memory_array[11411] <= 3'b000;
      memory_array[11412] <= 3'b000;
      memory_array[11413] <= 3'b000;
      memory_array[11414] <= 3'b000;
      memory_array[11415] <= 3'b000;
      memory_array[11416] <= 3'b000;
      memory_array[11417] <= 3'b000;
      memory_array[11418] <= 3'b110;
      memory_array[11419] <= 3'b000;
      memory_array[11420] <= 3'b101;
      memory_array[11421] <= 3'b000;
      memory_array[11422] <= 3'b000;
      memory_array[11423] <= 3'b101;
      memory_array[11424] <= 3'b000;
      memory_array[11425] <= 3'b101;
      memory_array[11426] <= 3'b000;
      memory_array[11427] <= 3'b101;
      memory_array[11428] <= 3'b101;
      memory_array[11429] <= 3'b101;
      memory_array[11430] <= 3'b000;
      memory_array[11431] <= 3'b000;
      memory_array[11432] <= 3'b000;
      memory_array[11433] <= 3'b000;
      memory_array[11434] <= 3'b101;
      memory_array[11435] <= 3'b111;
      memory_array[11436] <= 3'b111;
      memory_array[11437] <= 3'b111;
      memory_array[11438] <= 3'b111;
      memory_array[11439] <= 3'b000;
      memory_array[11440] <= 3'b101;
      memory_array[11441] <= 3'b101;
      memory_array[11442] <= 3'b101;
      memory_array[11443] <= 3'b101;
      memory_array[11444] <= 3'b101;
      memory_array[11445] <= 3'b101;
      memory_array[11446] <= 3'b101;
      memory_array[11447] <= 3'b101;
      memory_array[11448] <= 3'b101;
      memory_array[11449] <= 3'b101;
      memory_array[11450] <= 3'b101;
      memory_array[11451] <= 3'b101;
      memory_array[11452] <= 3'b101;
      memory_array[11453] <= 3'b000;
      memory_array[11454] <= 3'b000;
      memory_array[11455] <= 3'b000;
      memory_array[11456] <= 3'b000;
      memory_array[11457] <= 3'b000;
      memory_array[11458] <= 3'b101;
      memory_array[11459] <= 3'b000;
      memory_array[11460] <= 3'b101;
      memory_array[11461] <= 3'b101;
      memory_array[11462] <= 3'b101;
      memory_array[11463] <= 3'b101;
      memory_array[11464] <= 3'b101;
      memory_array[11465] <= 3'b101;
      memory_array[11466] <= 3'b111;
      memory_array[11467] <= 3'b101;
      memory_array[11468] <= 3'b111;
      memory_array[11469] <= 3'b101;
      memory_array[11470] <= 3'b101;
      memory_array[11471] <= 3'b101;
      memory_array[11472] <= 3'b101;
      memory_array[11473] <= 3'b101;
      memory_array[11474] <= 3'b111;
      memory_array[11475] <= 3'b111;
      memory_array[11476] <= 3'b111;
      memory_array[11477] <= 3'b111;
      memory_array[11478] <= 3'b111;
      memory_array[11479] <= 3'b111;
      memory_array[11480] <= 3'b101;
      memory_array[11481] <= 3'b111;
      memory_array[11482] <= 3'b111;
      memory_array[11483] <= 3'b101;
      memory_array[11484] <= 3'b111;
      memory_array[11485] <= 3'b111;
      memory_array[11486] <= 3'b101;
      memory_array[11487] <= 3'b000;
      memory_array[11488] <= 3'b101;
      memory_array[11489] <= 3'b111;
      memory_array[11490] <= 3'b111;
      memory_array[11491] <= 3'b111;
      memory_array[11492] <= 3'b000;
      memory_array[11493] <= 3'b101;
      memory_array[11494] <= 3'b110;
      memory_array[11495] <= 3'b111;
      memory_array[11496] <= 3'b111;
      memory_array[11497] <= 3'b111;
      memory_array[11498] <= 3'b111;
      memory_array[11499] <= 3'b111;
      memory_array[11500] <= 3'b111;
      memory_array[11501] <= 3'b111;
      memory_array[11502] <= 3'b101;
      memory_array[11503] <= 3'b111;
      memory_array[11504] <= 3'b101;
      memory_array[11505] <= 3'b111;
      memory_array[11506] <= 3'b111;
      memory_array[11507] <= 3'b000;
      memory_array[11508] <= 3'b000;
      memory_array[11509] <= 3'b000;
      memory_array[11510] <= 3'b000;
      memory_array[11511] <= 3'b000;
      memory_array[11512] <= 3'b000;
      memory_array[11513] <= 3'b000;
      memory_array[11514] <= 3'b101;
      memory_array[11515] <= 3'b101;
      memory_array[11516] <= 3'b101;
      memory_array[11517] <= 3'b111;
      memory_array[11518] <= 3'b111;
      memory_array[11519] <= 3'b101;
      memory_array[11520] <= 3'b101;
      memory_array[11521] <= 3'b110;
      memory_array[11522] <= 3'b101;
      memory_array[11523] <= 3'b101;
      memory_array[11524] <= 3'b101;
      memory_array[11525] <= 3'b101;
      memory_array[11526] <= 3'b101;
      memory_array[11527] <= 3'b101;
      memory_array[11528] <= 3'b101;
      memory_array[11529] <= 3'b101;
      memory_array[11530] <= 3'b101;
      memory_array[11531] <= 3'b101;
      memory_array[11532] <= 3'b101;
      memory_array[11533] <= 3'b110;
      memory_array[11534] <= 3'b101;
      memory_array[11535] <= 3'b101;
      memory_array[11536] <= 3'b101;
      memory_array[11537] <= 3'b101;
      memory_array[11538] <= 3'b101;
      memory_array[11539] <= 3'b101;
      memory_array[11540] <= 3'b101;
      memory_array[11541] <= 3'b101;
      memory_array[11542] <= 3'b110;
      memory_array[11543] <= 3'b110;
      memory_array[11544] <= 3'b110;
      memory_array[11545] <= 3'b110;
      memory_array[11546] <= 3'b110;
      memory_array[11547] <= 3'b110;
      memory_array[11548] <= 3'b110;
      memory_array[11549] <= 3'b110;
      memory_array[11550] <= 3'b110;
      memory_array[11551] <= 3'b101;
      memory_array[11552] <= 3'b101;
      memory_array[11553] <= 3'b101;
      memory_array[11554] <= 3'b101;
      memory_array[11555] <= 3'b101;
      memory_array[11556] <= 3'b101;
      memory_array[11557] <= 3'b101;
      memory_array[11558] <= 3'b101;
      memory_array[11559] <= 3'b101;
      memory_array[11560] <= 3'b000;
      memory_array[11561] <= 3'b111;
      memory_array[11562] <= 3'b111;
      memory_array[11563] <= 3'b111;
      memory_array[11564] <= 3'b111;
      memory_array[11565] <= 3'b101;
      memory_array[11566] <= 3'b000;
      memory_array[11567] <= 3'b101;
      memory_array[11568] <= 3'b000;
      memory_array[11569] <= 3'b000;
      memory_array[11570] <= 3'b101;
      memory_array[11571] <= 3'b000;
      memory_array[11572] <= 3'b000;
      memory_array[11573] <= 3'b000;
      memory_array[11574] <= 3'b101;
      memory_array[11575] <= 3'b000;
      memory_array[11576] <= 3'b101;
      memory_array[11577] <= 3'b000;
      memory_array[11578] <= 3'b000;
      memory_array[11579] <= 3'b101;
      memory_array[11580] <= 3'b000;
      memory_array[11581] <= 3'b000;
      memory_array[11582] <= 3'b000;
      memory_array[11583] <= 3'b110;
      memory_array[11584] <= 3'b110;
      memory_array[11585] <= 3'b000;
      memory_array[11586] <= 3'b000;
      memory_array[11587] <= 3'b000;
      memory_array[11588] <= 3'b110;
      memory_array[11589] <= 3'b000;
      memory_array[11590] <= 3'b000;
      memory_array[11591] <= 3'b101;
      memory_array[11592] <= 3'b000;
      memory_array[11593] <= 3'b110;
      memory_array[11594] <= 3'b110;
      memory_array[11595] <= 3'b000;
      memory_array[11596] <= 3'b000;
      memory_array[11597] <= 3'b000;
      memory_array[11598] <= 3'b110;
      memory_array[11599] <= 3'b110;
      memory_array[11600] <= 3'b101;
      memory_array[11601] <= 3'b101;
      memory_array[11602] <= 3'b101;
      memory_array[11603] <= 3'b101;
      memory_array[11604] <= 3'b101;
      memory_array[11605] <= 3'b101;
      memory_array[11606] <= 3'b101;
      memory_array[11607] <= 3'b101;
      memory_array[11608] <= 3'b101;
      memory_array[11609] <= 3'b000;
      memory_array[11610] <= 3'b000;
      memory_array[11611] <= 3'b110;
      memory_array[11612] <= 3'b110;
      memory_array[11613] <= 3'b000;
      memory_array[11614] <= 3'b000;
      memory_array[11615] <= 3'b110;
      memory_array[11616] <= 3'b110;
      memory_array[11617] <= 3'b110;
      memory_array[11618] <= 3'b000;
      memory_array[11619] <= 3'b000;
      memory_array[11620] <= 3'b110;
      memory_array[11621] <= 3'b110;
      memory_array[11622] <= 3'b000;
      memory_array[11623] <= 3'b101;
      memory_array[11624] <= 3'b000;
      memory_array[11625] <= 3'b000;
      memory_array[11626] <= 3'b000;
      memory_array[11627] <= 3'b101;
      memory_array[11628] <= 3'b101;
      memory_array[11629] <= 3'b101;
      memory_array[11630] <= 3'b000;
      memory_array[11631] <= 3'b000;
      memory_array[11632] <= 3'b101;
      memory_array[11633] <= 3'b000;
      memory_array[11634] <= 3'b000;
      memory_array[11635] <= 3'b111;
      memory_array[11636] <= 3'b111;
      memory_array[11637] <= 3'b111;
      memory_array[11638] <= 3'b111;
      memory_array[11639] <= 3'b000;
      memory_array[11640] <= 3'b101;
      memory_array[11641] <= 3'b101;
      memory_array[11642] <= 3'b101;
      memory_array[11643] <= 3'b101;
      memory_array[11644] <= 3'b101;
      memory_array[11645] <= 3'b101;
      memory_array[11646] <= 3'b101;
      memory_array[11647] <= 3'b101;
      memory_array[11648] <= 3'b101;
      memory_array[11649] <= 3'b101;
      memory_array[11650] <= 3'b101;
      memory_array[11651] <= 3'b101;
      memory_array[11652] <= 3'b000;
      memory_array[11653] <= 3'b000;
      memory_array[11654] <= 3'b000;
      memory_array[11655] <= 3'b000;
      memory_array[11656] <= 3'b000;
      memory_array[11657] <= 3'b000;
      memory_array[11658] <= 3'b000;
      memory_array[11659] <= 3'b000;
      memory_array[11660] <= 3'b000;
      memory_array[11661] <= 3'b101;
      memory_array[11662] <= 3'b101;
      memory_array[11663] <= 3'b101;
      memory_array[11664] <= 3'b101;
      memory_array[11665] <= 3'b101;
      memory_array[11666] <= 3'b111;
      memory_array[11667] <= 3'b101;
      memory_array[11668] <= 3'b101;
      memory_array[11669] <= 3'b000;
      memory_array[11670] <= 3'b000;
      memory_array[11671] <= 3'b111;
      memory_array[11672] <= 3'b101;
      memory_array[11673] <= 3'b111;
      memory_array[11674] <= 3'b101;
      memory_array[11675] <= 3'b111;
      memory_array[11676] <= 3'b111;
      memory_array[11677] <= 3'b111;
      memory_array[11678] <= 3'b111;
      memory_array[11679] <= 3'b111;
      memory_array[11680] <= 3'b101;
      memory_array[11681] <= 3'b111;
      memory_array[11682] <= 3'b111;
      memory_array[11683] <= 3'b101;
      memory_array[11684] <= 3'b111;
      memory_array[11685] <= 3'b111;
      memory_array[11686] <= 3'b101;
      memory_array[11687] <= 3'b000;
      memory_array[11688] <= 3'b000;
      memory_array[11689] <= 3'b000;
      memory_array[11690] <= 3'b101;
      memory_array[11691] <= 3'b111;
      memory_array[11692] <= 3'b101;
      memory_array[11693] <= 3'b101;
      memory_array[11694] <= 3'b000;
      memory_array[11695] <= 3'b110;
      memory_array[11696] <= 3'b111;
      memory_array[11697] <= 3'b111;
      memory_array[11698] <= 3'b111;
      memory_array[11699] <= 3'b111;
      memory_array[11700] <= 3'b111;
      memory_array[11701] <= 3'b111;
      memory_array[11702] <= 3'b101;
      memory_array[11703] <= 3'b111;
      memory_array[11704] <= 3'b000;
      memory_array[11705] <= 3'b101;
      memory_array[11706] <= 3'b111;
      memory_array[11707] <= 3'b101;
      memory_array[11708] <= 3'b000;
      memory_array[11709] <= 3'b000;
      memory_array[11710] <= 3'b000;
      memory_array[11711] <= 3'b101;
      memory_array[11712] <= 3'b000;
      memory_array[11713] <= 3'b000;
      memory_array[11714] <= 3'b000;
      memory_array[11715] <= 3'b000;
      memory_array[11716] <= 3'b101;
      memory_array[11717] <= 3'b111;
      memory_array[11718] <= 3'b111;
      memory_array[11719] <= 3'b111;
      memory_array[11720] <= 3'b101;
      memory_array[11721] <= 3'b110;
      memory_array[11722] <= 3'b101;
      memory_array[11723] <= 3'b101;
      memory_array[11724] <= 3'b101;
      memory_array[11725] <= 3'b101;
      memory_array[11726] <= 3'b101;
      memory_array[11727] <= 3'b101;
      memory_array[11728] <= 3'b101;
      memory_array[11729] <= 3'b101;
      memory_array[11730] <= 3'b101;
      memory_array[11731] <= 3'b101;
      memory_array[11732] <= 3'b110;
      memory_array[11733] <= 3'b110;
      memory_array[11734] <= 3'b110;
      memory_array[11735] <= 3'b110;
      memory_array[11736] <= 3'b110;
      memory_array[11737] <= 3'b110;
      memory_array[11738] <= 3'b000;
      memory_array[11739] <= 3'b000;
      memory_array[11740] <= 3'b000;
      memory_array[11741] <= 3'b110;
      memory_array[11742] <= 3'b110;
      memory_array[11743] <= 3'b101;
      memory_array[11744] <= 3'b101;
      memory_array[11745] <= 3'b110;
      memory_array[11746] <= 3'b110;
      memory_array[11747] <= 3'b110;
      memory_array[11748] <= 3'b000;
      memory_array[11749] <= 3'b000;
      memory_array[11750] <= 3'b110;
      memory_array[11751] <= 3'b110;
      memory_array[11752] <= 3'b000;
      memory_array[11753] <= 3'b000;
      memory_array[11754] <= 3'b101;
      memory_array[11755] <= 3'b101;
      memory_array[11756] <= 3'b101;
      memory_array[11757] <= 3'b101;
      memory_array[11758] <= 3'b101;
      memory_array[11759] <= 3'b101;
      memory_array[11760] <= 3'b000;
      memory_array[11761] <= 3'b111;
      memory_array[11762] <= 3'b111;
      memory_array[11763] <= 3'b111;
      memory_array[11764] <= 3'b111;
      memory_array[11765] <= 3'b000;
      memory_array[11766] <= 3'b000;
      memory_array[11767] <= 3'b101;
      memory_array[11768] <= 3'b000;
      memory_array[11769] <= 3'b000;
      memory_array[11770] <= 3'b101;
      memory_array[11771] <= 3'b101;
      memory_array[11772] <= 3'b000;
      memory_array[11773] <= 3'b000;
      memory_array[11774] <= 3'b000;
      memory_array[11775] <= 3'b000;
      memory_array[11776] <= 3'b101;
      memory_array[11777] <= 3'b000;
      memory_array[11778] <= 3'b000;
      memory_array[11779] <= 3'b000;
      memory_array[11780] <= 3'b000;
      memory_array[11781] <= 3'b110;
      memory_array[11782] <= 3'b110;
      memory_array[11783] <= 3'b000;
      memory_array[11784] <= 3'b000;
      memory_array[11785] <= 3'b110;
      memory_array[11786] <= 3'b000;
      memory_array[11787] <= 3'b110;
      memory_array[11788] <= 3'b000;
      memory_array[11789] <= 3'b000;
      memory_array[11790] <= 3'b000;
      memory_array[11791] <= 3'b101;
      memory_array[11792] <= 3'b101;
      memory_array[11793] <= 3'b101;
      memory_array[11794] <= 3'b101;
      memory_array[11795] <= 3'b101;
      memory_array[11796] <= 3'b101;
      memory_array[11797] <= 3'b101;
      memory_array[11798] <= 3'b101;
      memory_array[11799] <= 3'b101;
      memory_array[11800] <= 3'b101;
      memory_array[11801] <= 3'b101;
      memory_array[11802] <= 3'b101;
      memory_array[11803] <= 3'b101;
      memory_array[11804] <= 3'b101;
      memory_array[11805] <= 3'b101;
      memory_array[11806] <= 3'b101;
      memory_array[11807] <= 3'b101;
      memory_array[11808] <= 3'b101;
      memory_array[11809] <= 3'b000;
      memory_array[11810] <= 3'b000;
      memory_array[11811] <= 3'b110;
      memory_array[11812] <= 3'b111;
      memory_array[11813] <= 3'b000;
      memory_array[11814] <= 3'b000;
      memory_array[11815] <= 3'b101;
      memory_array[11816] <= 3'b110;
      memory_array[11817] <= 3'b000;
      memory_array[11818] <= 3'b101;
      memory_array[11819] <= 3'b101;
      memory_array[11820] <= 3'b000;
      memory_array[11821] <= 3'b110;
      memory_array[11822] <= 3'b101;
      memory_array[11823] <= 3'b000;
      memory_array[11824] <= 3'b000;
      memory_array[11825] <= 3'b000;
      memory_array[11826] <= 3'b110;
      memory_array[11827] <= 3'b000;
      memory_array[11828] <= 3'b000;
      memory_array[11829] <= 3'b101;
      memory_array[11830] <= 3'b101;
      memory_array[11831] <= 3'b110;
      memory_array[11832] <= 3'b110;
      memory_array[11833] <= 3'b000;
      memory_array[11834] <= 3'b000;
      memory_array[11835] <= 3'b000;
      memory_array[11836] <= 3'b111;
      memory_array[11837] <= 3'b111;
      memory_array[11838] <= 3'b111;
      memory_array[11839] <= 3'b101;
      memory_array[11840] <= 3'b000;
      memory_array[11841] <= 3'b101;
      memory_array[11842] <= 3'b101;
      memory_array[11843] <= 3'b000;
      memory_array[11844] <= 3'b000;
      memory_array[11845] <= 3'b101;
      memory_array[11846] <= 3'b101;
      memory_array[11847] <= 3'b101;
      memory_array[11848] <= 3'b000;
      memory_array[11849] <= 3'b000;
      memory_array[11850] <= 3'b000;
      memory_array[11851] <= 3'b000;
      memory_array[11852] <= 3'b000;
      memory_array[11853] <= 3'b000;
      memory_array[11854] <= 3'b000;
      memory_array[11855] <= 3'b000;
      memory_array[11856] <= 3'b000;
      memory_array[11857] <= 3'b101;
      memory_array[11858] <= 3'b000;
      memory_array[11859] <= 3'b000;
      memory_array[11860] <= 3'b101;
      memory_array[11861] <= 3'b101;
      memory_array[11862] <= 3'b101;
      memory_array[11863] <= 3'b000;
      memory_array[11864] <= 3'b000;
      memory_array[11865] <= 3'b101;
      memory_array[11866] <= 3'b111;
      memory_array[11867] <= 3'b101;
      memory_array[11868] <= 3'b000;
      memory_array[11869] <= 3'b000;
      memory_array[11870] <= 3'b101;
      memory_array[11871] <= 3'b000;
      memory_array[11872] <= 3'b111;
      memory_array[11873] <= 3'b111;
      memory_array[11874] <= 3'b111;
      memory_array[11875] <= 3'b111;
      memory_array[11876] <= 3'b111;
      memory_array[11877] <= 3'b111;
      memory_array[11878] <= 3'b111;
      memory_array[11879] <= 3'b101;
      memory_array[11880] <= 3'b000;
      memory_array[11881] <= 3'b111;
      memory_array[11882] <= 3'b111;
      memory_array[11883] <= 3'b111;
      memory_array[11884] <= 3'b111;
      memory_array[11885] <= 3'b111;
      memory_array[11886] <= 3'b101;
      memory_array[11887] <= 3'b101;
      memory_array[11888] <= 3'b000;
      memory_array[11889] <= 3'b000;
      memory_array[11890] <= 3'b101;
      memory_array[11891] <= 3'b000;
      memory_array[11892] <= 3'b110;
      memory_array[11893] <= 3'b000;
      memory_array[11894] <= 3'b000;
      memory_array[11895] <= 3'b110;
      memory_array[11896] <= 3'b110;
      memory_array[11897] <= 3'b111;
      memory_array[11898] <= 3'b111;
      memory_array[11899] <= 3'b111;
      memory_array[11900] <= 3'b111;
      memory_array[11901] <= 3'b111;
      memory_array[11902] <= 3'b101;
      memory_array[11903] <= 3'b000;
      memory_array[11904] <= 3'b000;
      memory_array[11905] <= 3'b111;
      memory_array[11906] <= 3'b111;
      memory_array[11907] <= 3'b000;
      memory_array[11908] <= 3'b000;
      memory_array[11909] <= 3'b000;
      memory_array[11910] <= 3'b101;
      memory_array[11911] <= 3'b101;
      memory_array[11912] <= 3'b000;
      memory_array[11913] <= 3'b000;
      memory_array[11914] <= 3'b000;
      memory_array[11915] <= 3'b000;
      memory_array[11916] <= 3'b000;
      memory_array[11917] <= 3'b000;
      memory_array[11918] <= 3'b111;
      memory_array[11919] <= 3'b111;
      memory_array[11920] <= 3'b101;
      memory_array[11921] <= 3'b110;
      memory_array[11922] <= 3'b101;
      memory_array[11923] <= 3'b000;
      memory_array[11924] <= 3'b000;
      memory_array[11925] <= 3'b101;
      memory_array[11926] <= 3'b101;
      memory_array[11927] <= 3'b101;
      memory_array[11928] <= 3'b000;
      memory_array[11929] <= 3'b000;
      memory_array[11930] <= 3'b101;
      memory_array[11931] <= 3'b101;
      memory_array[11932] <= 3'b101;
      memory_array[11933] <= 3'b000;
      memory_array[11934] <= 3'b110;
      memory_array[11935] <= 3'b101;
      memory_array[11936] <= 3'b101;
      memory_array[11937] <= 3'b101;
      memory_array[11938] <= 3'b000;
      memory_array[11939] <= 3'b000;
      memory_array[11940] <= 3'b110;
      memory_array[11941] <= 3'b110;
      memory_array[11942] <= 3'b110;
      memory_array[11943] <= 3'b000;
      memory_array[11944] <= 3'b000;
      memory_array[11945] <= 3'b110;
      memory_array[11946] <= 3'b101;
      memory_array[11947] <= 3'b101;
      memory_array[11948] <= 3'b000;
      memory_array[11949] <= 3'b000;
      memory_array[11950] <= 3'b101;
      memory_array[11951] <= 3'b101;
      memory_array[11952] <= 3'b101;
      memory_array[11953] <= 3'b000;
      memory_array[11954] <= 3'b000;
      memory_array[11955] <= 3'b101;
      memory_array[11956] <= 3'b101;
      memory_array[11957] <= 3'b101;
      memory_array[11958] <= 3'b000;
      memory_array[11959] <= 3'b000;
      memory_array[11960] <= 3'b101;
      memory_array[11961] <= 3'b111;
      memory_array[11962] <= 3'b111;
      memory_array[11963] <= 3'b111;
      memory_array[11964] <= 3'b000;
      memory_array[11965] <= 3'b110;
      memory_array[11966] <= 3'b110;
      memory_array[11967] <= 3'b000;
      memory_array[11968] <= 3'b000;
      memory_array[11969] <= 3'b101;
      memory_array[11970] <= 3'b101;
      memory_array[11971] <= 3'b000;
      memory_array[11972] <= 3'b110;
      memory_array[11973] <= 3'b000;
      memory_array[11974] <= 3'b000;
      memory_array[11975] <= 3'b110;
      memory_array[11976] <= 3'b000;
      memory_array[11977] <= 3'b000;
      memory_array[11978] <= 3'b000;
      memory_array[11979] <= 3'b000;
      memory_array[11980] <= 3'b101;
      memory_array[11981] <= 3'b101;
      memory_array[11982] <= 3'b110;
      memory_array[11983] <= 3'b000;
      memory_array[11984] <= 3'b101;
      memory_array[11985] <= 3'b000;
      memory_array[11986] <= 3'b000;
      memory_array[11987] <= 3'b000;
      memory_array[11988] <= 3'b000;
      memory_array[11989] <= 3'b000;
      memory_array[11990] <= 3'b000;
      memory_array[11991] <= 3'b101;
      memory_array[11992] <= 3'b101;
      memory_array[11993] <= 3'b101;
      memory_array[11994] <= 3'b101;
      memory_array[11995] <= 3'b101;
      memory_array[11996] <= 3'b101;
      memory_array[11997] <= 3'b101;
      memory_array[11998] <= 3'b101;
      memory_array[11999] <= 3'b101;
      memory_array[12000] <= 3'b000;
      memory_array[12001] <= 3'b000;
      memory_array[12002] <= 3'b000;
      memory_array[12003] <= 3'b110;
      memory_array[12004] <= 3'b110;
      memory_array[12005] <= 3'b000;
      memory_array[12006] <= 3'b000;
      memory_array[12007] <= 3'b000;
      memory_array[12008] <= 3'b101;
      memory_array[12009] <= 3'b000;
      memory_array[12010] <= 3'b000;
      memory_array[12011] <= 3'b101;
      memory_array[12012] <= 3'b000;
      memory_array[12013] <= 3'b111;
      memory_array[12014] <= 3'b101;
      memory_array[12015] <= 3'b000;
      memory_array[12016] <= 3'b101;
      memory_array[12017] <= 3'b000;
      memory_array[12018] <= 3'b101;
      memory_array[12019] <= 3'b000;
      memory_array[12020] <= 3'b101;
      memory_array[12021] <= 3'b000;
      memory_array[12022] <= 3'b000;
      memory_array[12023] <= 3'b000;
      memory_array[12024] <= 3'b000;
      memory_array[12025] <= 3'b101;
      memory_array[12026] <= 3'b101;
      memory_array[12027] <= 3'b000;
      memory_array[12028] <= 3'b000;
      memory_array[12029] <= 3'b000;
      memory_array[12030] <= 3'b101;
      memory_array[12031] <= 3'b000;
      memory_array[12032] <= 3'b000;
      memory_array[12033] <= 3'b110;
      memory_array[12034] <= 3'b110;
      memory_array[12035] <= 3'b000;
      memory_array[12036] <= 3'b111;
      memory_array[12037] <= 3'b111;
      memory_array[12038] <= 3'b111;
      memory_array[12039] <= 3'b111;
      memory_array[12040] <= 3'b000;
      memory_array[12041] <= 3'b000;
      memory_array[12042] <= 3'b110;
      memory_array[12043] <= 3'b110;
      memory_array[12044] <= 3'b101;
      memory_array[12045] <= 3'b000;
      memory_array[12046] <= 3'b000;
      memory_array[12047] <= 3'b000;
      memory_array[12048] <= 3'b000;
      memory_array[12049] <= 3'b000;
      memory_array[12050] <= 3'b000;
      memory_array[12051] <= 3'b000;
      memory_array[12052] <= 3'b000;
      memory_array[12053] <= 3'b000;
      memory_array[12054] <= 3'b000;
      memory_array[12055] <= 3'b000;
      memory_array[12056] <= 3'b000;
      memory_array[12057] <= 3'b000;
      memory_array[12058] <= 3'b000;
      memory_array[12059] <= 3'b101;
      memory_array[12060] <= 3'b000;
      memory_array[12061] <= 3'b000;
      memory_array[12062] <= 3'b000;
      memory_array[12063] <= 3'b101;
      memory_array[12064] <= 3'b101;
      memory_array[12065] <= 3'b000;
      memory_array[12066] <= 3'b111;
      memory_array[12067] <= 3'b000;
      memory_array[12068] <= 3'b101;
      memory_array[12069] <= 3'b000;
      memory_array[12070] <= 3'b000;
      memory_array[12071] <= 3'b000;
      memory_array[12072] <= 3'b000;
      memory_array[12073] <= 3'b101;
      memory_array[12074] <= 3'b111;
      memory_array[12075] <= 3'b111;
      memory_array[12076] <= 3'b111;
      memory_array[12077] <= 3'b101;
      memory_array[12078] <= 3'b101;
      memory_array[12079] <= 3'b000;
      memory_array[12080] <= 3'b000;
      memory_array[12081] <= 3'b111;
      memory_array[12082] <= 3'b000;
      memory_array[12083] <= 3'b000;
      memory_array[12084] <= 3'b101;
      memory_array[12085] <= 3'b000;
      memory_array[12086] <= 3'b111;
      memory_array[12087] <= 3'b111;
      memory_array[12088] <= 3'b111;
      memory_array[12089] <= 3'b111;
      memory_array[12090] <= 3'b111;
      memory_array[12091] <= 3'b000;
      memory_array[12092] <= 3'b000;
      memory_array[12093] <= 3'b110;
      memory_array[12094] <= 3'b110;
      memory_array[12095] <= 3'b000;
      memory_array[12096] <= 3'b000;
      memory_array[12097] <= 3'b000;
      memory_array[12098] <= 3'b111;
      memory_array[12099] <= 3'b111;
      memory_array[12100] <= 3'b111;
      memory_array[12101] <= 3'b000;
      memory_array[12102] <= 3'b000;
      memory_array[12103] <= 3'b101;
      memory_array[12104] <= 3'b101;
      memory_array[12105] <= 3'b000;
      memory_array[12106] <= 3'b000;
      memory_array[12107] <= 3'b000;
      memory_array[12108] <= 3'b000;
      memory_array[12109] <= 3'b101;
      memory_array[12110] <= 3'b000;
      memory_array[12111] <= 3'b000;
      memory_array[12112] <= 3'b000;
      memory_array[12113] <= 3'b000;
      memory_array[12114] <= 3'b101;
      memory_array[12115] <= 3'b000;
      memory_array[12116] <= 3'b000;
      memory_array[12117] <= 3'b000;
      memory_array[12118] <= 3'b000;
      memory_array[12119] <= 3'b000;
      memory_array[12120] <= 3'b101;
      memory_array[12121] <= 3'b110;
      memory_array[12122] <= 3'b000;
      memory_array[12123] <= 3'b101;
      memory_array[12124] <= 3'b101;
      memory_array[12125] <= 3'b000;
      memory_array[12126] <= 3'b000;
      memory_array[12127] <= 3'b000;
      memory_array[12128] <= 3'b101;
      memory_array[12129] <= 3'b101;
      memory_array[12130] <= 3'b000;
      memory_array[12131] <= 3'b000;
      memory_array[12132] <= 3'b000;
      memory_array[12133] <= 3'b101;
      memory_array[12134] <= 3'b101;
      memory_array[12135] <= 3'b000;
      memory_array[12136] <= 3'b000;
      memory_array[12137] <= 3'b000;
      memory_array[12138] <= 3'b101;
      memory_array[12139] <= 3'b101;
      memory_array[12140] <= 3'b000;
      memory_array[12141] <= 3'b000;
      memory_array[12142] <= 3'b000;
      memory_array[12143] <= 3'b101;
      memory_array[12144] <= 3'b101;
      memory_array[12145] <= 3'b000;
      memory_array[12146] <= 3'b110;
      memory_array[12147] <= 3'b000;
      memory_array[12148] <= 3'b101;
      memory_array[12149] <= 3'b101;
      memory_array[12150] <= 3'b000;
      memory_array[12151] <= 3'b000;
      memory_array[12152] <= 3'b110;
      memory_array[12153] <= 3'b101;
      memory_array[12154] <= 3'b101;
      memory_array[12155] <= 3'b000;
      memory_array[12156] <= 3'b000;
      memory_array[12157] <= 3'b000;
      memory_array[12158] <= 3'b101;
      memory_array[12159] <= 3'b000;
      memory_array[12160] <= 3'b111;
      memory_array[12161] <= 3'b111;
      memory_array[12162] <= 3'b111;
      memory_array[12163] <= 3'b111;
      memory_array[12164] <= 3'b000;
      memory_array[12165] <= 3'b000;
      memory_array[12166] <= 3'b000;
      memory_array[12167] <= 3'b000;
      memory_array[12168] <= 3'b000;
      memory_array[12169] <= 3'b101;
      memory_array[12170] <= 3'b000;
      memory_array[12171] <= 3'b000;
      memory_array[12172] <= 3'b000;
      memory_array[12173] <= 3'b101;
      memory_array[12174] <= 3'b101;
      memory_array[12175] <= 3'b000;
      memory_array[12176] <= 3'b000;
      memory_array[12177] <= 3'b101;
      memory_array[12178] <= 3'b000;
      memory_array[12179] <= 3'b101;
      memory_array[12180] <= 3'b000;
      memory_array[12181] <= 3'b101;
      memory_array[12182] <= 3'b000;
      memory_array[12183] <= 3'b101;
      memory_array[12184] <= 3'b000;
      memory_array[12185] <= 3'b101;
      memory_array[12186] <= 3'b111;
      memory_array[12187] <= 3'b101;
      memory_array[12188] <= 3'b101;
      memory_array[12189] <= 3'b000;
      memory_array[12190] <= 3'b000;
      memory_array[12191] <= 3'b101;
      memory_array[12192] <= 3'b000;
      memory_array[12193] <= 3'b110;
      memory_array[12194] <= 3'b110;
      memory_array[12195] <= 3'b000;
      memory_array[12196] <= 3'b000;
      memory_array[12197] <= 3'b000;
      memory_array[12198] <= 3'b110;
      memory_array[12199] <= 3'b110;
      memory_array[12200] <= 3'b101;
      memory_array[12201] <= 3'b110;
      memory_array[12202] <= 3'b110;
      memory_array[12203] <= 3'b000;
      memory_array[12204] <= 3'b000;
      memory_array[12205] <= 3'b110;
      memory_array[12206] <= 3'b110;
      memory_array[12207] <= 3'b101;
      memory_array[12208] <= 3'b101;
      memory_array[12209] <= 3'b000;
      memory_array[12210] <= 3'b000;
      memory_array[12211] <= 3'b000;
      memory_array[12212] <= 3'b101;
      memory_array[12213] <= 3'b000;
      memory_array[12214] <= 3'b000;
      memory_array[12215] <= 3'b101;
      memory_array[12216] <= 3'b110;
      memory_array[12217] <= 3'b000;
      memory_array[12218] <= 3'b000;
      memory_array[12219] <= 3'b000;
      memory_array[12220] <= 3'b000;
      memory_array[12221] <= 3'b101;
      memory_array[12222] <= 3'b000;
      memory_array[12223] <= 3'b000;
      memory_array[12224] <= 3'b101;
      memory_array[12225] <= 3'b101;
      memory_array[12226] <= 3'b101;
      memory_array[12227] <= 3'b000;
      memory_array[12228] <= 3'b000;
      memory_array[12229] <= 3'b000;
      memory_array[12230] <= 3'b000;
      memory_array[12231] <= 3'b101;
      memory_array[12232] <= 3'b000;
      memory_array[12233] <= 3'b000;
      memory_array[12234] <= 3'b000;
      memory_array[12235] <= 3'b110;
      memory_array[12236] <= 3'b111;
      memory_array[12237] <= 3'b111;
      memory_array[12238] <= 3'b111;
      memory_array[12239] <= 3'b111;
      memory_array[12240] <= 3'b101;
      memory_array[12241] <= 3'b000;
      memory_array[12242] <= 3'b101;
      memory_array[12243] <= 3'b000;
      memory_array[12244] <= 3'b000;
      memory_array[12245] <= 3'b000;
      memory_array[12246] <= 3'b000;
      memory_array[12247] <= 3'b000;
      memory_array[12248] <= 3'b000;
      memory_array[12249] <= 3'b000;
      memory_array[12250] <= 3'b000;
      memory_array[12251] <= 3'b000;
      memory_array[12252] <= 3'b000;
      memory_array[12253] <= 3'b000;
      memory_array[12254] <= 3'b000;
      memory_array[12255] <= 3'b000;
      memory_array[12256] <= 3'b101;
      memory_array[12257] <= 3'b000;
      memory_array[12258] <= 3'b000;
      memory_array[12259] <= 3'b000;
      memory_array[12260] <= 3'b101;
      memory_array[12261] <= 3'b101;
      memory_array[12262] <= 3'b101;
      memory_array[12263] <= 3'b000;
      memory_array[12264] <= 3'b000;
      memory_array[12265] <= 3'b000;
      memory_array[12266] <= 3'b000;
      memory_array[12267] <= 3'b101;
      memory_array[12268] <= 3'b101;
      memory_array[12269] <= 3'b000;
      memory_array[12270] <= 3'b101;
      memory_array[12271] <= 3'b101;
      memory_array[12272] <= 3'b101;
      memory_array[12273] <= 3'b000;
      memory_array[12274] <= 3'b000;
      memory_array[12275] <= 3'b000;
      memory_array[12276] <= 3'b101;
      memory_array[12277] <= 3'b101;
      memory_array[12278] <= 3'b101;
      memory_array[12279] <= 3'b000;
      memory_array[12280] <= 3'b000;
      memory_array[12281] <= 3'b101;
      memory_array[12282] <= 3'b000;
      memory_array[12283] <= 3'b101;
      memory_array[12284] <= 3'b000;
      memory_array[12285] <= 3'b101;
      memory_array[12286] <= 3'b000;
      memory_array[12287] <= 3'b000;
      memory_array[12288] <= 3'b000;
      memory_array[12289] <= 3'b000;
      memory_array[12290] <= 3'b101;
      memory_array[12291] <= 3'b000;
      memory_array[12292] <= 3'b111;
      memory_array[12293] <= 3'b111;
      memory_array[12294] <= 3'b111;
      memory_array[12295] <= 3'b101;
      memory_array[12296] <= 3'b101;
      memory_array[12297] <= 3'b000;
      memory_array[12298] <= 3'b000;
      memory_array[12299] <= 3'b000;
      memory_array[12300] <= 3'b101;
      memory_array[12301] <= 3'b101;
      memory_array[12302] <= 3'b101;
      memory_array[12303] <= 3'b000;
      memory_array[12304] <= 3'b000;
      memory_array[12305] <= 3'b101;
      memory_array[12306] <= 3'b101;
      memory_array[12307] <= 3'b000;
      memory_array[12308] <= 3'b000;
      memory_array[12309] <= 3'b000;
      memory_array[12310] <= 3'b000;
      memory_array[12311] <= 3'b000;
      memory_array[12312] <= 3'b101;
      memory_array[12313] <= 3'b000;
      memory_array[12314] <= 3'b000;
      memory_array[12315] <= 3'b101;
      memory_array[12316] <= 3'b101;
      memory_array[12317] <= 3'b000;
      memory_array[12318] <= 3'b000;
      memory_array[12319] <= 3'b000;
      memory_array[12320] <= 3'b000;
      memory_array[12321] <= 3'b000;
      memory_array[12322] <= 3'b101;
      memory_array[12323] <= 3'b000;
      memory_array[12324] <= 3'b000;
      memory_array[12325] <= 3'b101;
      memory_array[12326] <= 3'b101;
      memory_array[12327] <= 3'b101;
      memory_array[12328] <= 3'b000;
      memory_array[12329] <= 3'b000;
      memory_array[12330] <= 3'b101;
      memory_array[12331] <= 3'b101;
      memory_array[12332] <= 3'b101;
      memory_array[12333] <= 3'b000;
      memory_array[12334] <= 3'b000;
      memory_array[12335] <= 3'b101;
      memory_array[12336] <= 3'b000;
      memory_array[12337] <= 3'b000;
      memory_array[12338] <= 3'b000;
      memory_array[12339] <= 3'b000;
      memory_array[12340] <= 3'b000;
      memory_array[12341] <= 3'b000;
      memory_array[12342] <= 3'b000;
      memory_array[12343] <= 3'b000;
      memory_array[12344] <= 3'b000;
      memory_array[12345] <= 3'b000;
      memory_array[12346] <= 3'b000;
      memory_array[12347] <= 3'b110;
      memory_array[12348] <= 3'b110;
      memory_array[12349] <= 3'b110;
      memory_array[12350] <= 3'b101;
      memory_array[12351] <= 3'b110;
      memory_array[12352] <= 3'b101;
      memory_array[12353] <= 3'b000;
      memory_array[12354] <= 3'b000;
      memory_array[12355] <= 3'b101;
      memory_array[12356] <= 3'b101;
      memory_array[12357] <= 3'b101;
      memory_array[12358] <= 3'b000;
      memory_array[12359] <= 3'b101;
      memory_array[12360] <= 3'b111;
      memory_array[12361] <= 3'b111;
      memory_array[12362] <= 3'b111;
      memory_array[12363] <= 3'b111;
      memory_array[12364] <= 3'b000;
      memory_array[12365] <= 3'b110;
      memory_array[12366] <= 3'b110;
      memory_array[12367] <= 3'b101;
      memory_array[12368] <= 3'b101;
      memory_array[12369] <= 3'b000;
      memory_array[12370] <= 3'b000;
      memory_array[12371] <= 3'b000;
      memory_array[12372] <= 3'b101;
      memory_array[12373] <= 3'b101;
      memory_array[12374] <= 3'b101;
      memory_array[12375] <= 3'b101;
      memory_array[12376] <= 3'b110;
      memory_array[12377] <= 3'b101;
      memory_array[12378] <= 3'b101;
      memory_array[12379] <= 3'b000;
      memory_array[12380] <= 3'b000;
      memory_array[12381] <= 3'b110;
      memory_array[12382] <= 3'b110;
      memory_array[12383] <= 3'b000;
      memory_array[12384] <= 3'b101;
      memory_array[12385] <= 3'b000;
      memory_array[12386] <= 3'b000;
      memory_array[12387] <= 3'b000;
      memory_array[12388] <= 3'b000;
      memory_array[12389] <= 3'b000;
      memory_array[12390] <= 3'b000;
      memory_array[12391] <= 3'b101;
      memory_array[12392] <= 3'b110;
      memory_array[12393] <= 3'b000;
      memory_array[12394] <= 3'b000;
      memory_array[12395] <= 3'b110;
      memory_array[12396] <= 3'b110;
      memory_array[12397] <= 3'b110;
      memory_array[12398] <= 3'b000;
      memory_array[12399] <= 3'b101;
      memory_array[12400] <= 3'b101;
      memory_array[12401] <= 3'b101;
      memory_array[12402] <= 3'b110;
      memory_array[12403] <= 3'b101;
      memory_array[12404] <= 3'b101;
      memory_array[12405] <= 3'b110;
      memory_array[12406] <= 3'b101;
      memory_array[12407] <= 3'b101;
      memory_array[12408] <= 3'b101;
      memory_array[12409] <= 3'b000;
      memory_array[12410] <= 3'b000;
      memory_array[12411] <= 3'b110;
      memory_array[12412] <= 3'b111;
      memory_array[12413] <= 3'b000;
      memory_array[12414] <= 3'b000;
      memory_array[12415] <= 3'b101;
      memory_array[12416] <= 3'b000;
      memory_array[12417] <= 3'b000;
      memory_array[12418] <= 3'b000;
      memory_array[12419] <= 3'b000;
      memory_array[12420] <= 3'b000;
      memory_array[12421] <= 3'b000;
      memory_array[12422] <= 3'b000;
      memory_array[12423] <= 3'b000;
      memory_array[12424] <= 3'b000;
      memory_array[12425] <= 3'b101;
      memory_array[12426] <= 3'b000;
      memory_array[12427] <= 3'b101;
      memory_array[12428] <= 3'b000;
      memory_array[12429] <= 3'b000;
      memory_array[12430] <= 3'b110;
      memory_array[12431] <= 3'b000;
      memory_array[12432] <= 3'b000;
      memory_array[12433] <= 3'b000;
      memory_array[12434] <= 3'b000;
      memory_array[12435] <= 3'b000;
      memory_array[12436] <= 3'b000;
      memory_array[12437] <= 3'b111;
      memory_array[12438] <= 3'b111;
      memory_array[12439] <= 3'b111;
      memory_array[12440] <= 3'b111;
      memory_array[12441] <= 3'b101;
      memory_array[12442] <= 3'b000;
      memory_array[12443] <= 3'b000;
      memory_array[12444] <= 3'b000;
      memory_array[12445] <= 3'b000;
      memory_array[12446] <= 3'b000;
      memory_array[12447] <= 3'b000;
      memory_array[12448] <= 3'b000;
      memory_array[12449] <= 3'b000;
      memory_array[12450] <= 3'b000;
      memory_array[12451] <= 3'b000;
      memory_array[12452] <= 3'b000;
      memory_array[12453] <= 3'b000;
      memory_array[12454] <= 3'b000;
      memory_array[12455] <= 3'b101;
      memory_array[12456] <= 3'b101;
      memory_array[12457] <= 3'b000;
      memory_array[12458] <= 3'b000;
      memory_array[12459] <= 3'b000;
      memory_array[12460] <= 3'b000;
      memory_array[12461] <= 3'b000;
      memory_array[12462] <= 3'b101;
      memory_array[12463] <= 3'b000;
      memory_array[12464] <= 3'b000;
      memory_array[12465] <= 3'b000;
      memory_array[12466] <= 3'b101;
      memory_array[12467] <= 3'b101;
      memory_array[12468] <= 3'b101;
      memory_array[12469] <= 3'b111;
      memory_array[12470] <= 3'b101;
      memory_array[12471] <= 3'b101;
      memory_array[12472] <= 3'b101;
      memory_array[12473] <= 3'b000;
      memory_array[12474] <= 3'b000;
      memory_array[12475] <= 3'b101;
      memory_array[12476] <= 3'b101;
      memory_array[12477] <= 3'b101;
      memory_array[12478] <= 3'b000;
      memory_array[12479] <= 3'b000;
      memory_array[12480] <= 3'b101;
      memory_array[12481] <= 3'b101;
      memory_array[12482] <= 3'b111;
      memory_array[12483] <= 3'b000;
      memory_array[12484] <= 3'b101;
      memory_array[12485] <= 3'b000;
      memory_array[12486] <= 3'b000;
      memory_array[12487] <= 3'b101;
      memory_array[12488] <= 3'b000;
      memory_array[12489] <= 3'b000;
      memory_array[12490] <= 3'b101;
      memory_array[12491] <= 3'b101;
      memory_array[12492] <= 3'b111;
      memory_array[12493] <= 3'b111;
      memory_array[12494] <= 3'b101;
      memory_array[12495] <= 3'b101;
      memory_array[12496] <= 3'b111;
      memory_array[12497] <= 3'b000;
      memory_array[12498] <= 3'b000;
      memory_array[12499] <= 3'b000;
      memory_array[12500] <= 3'b101;
      memory_array[12501] <= 3'b101;
      memory_array[12502] <= 3'b000;
      memory_array[12503] <= 3'b000;
      memory_array[12504] <= 3'b000;
      memory_array[12505] <= 3'b111;
      memory_array[12506] <= 3'b111;
      memory_array[12507] <= 3'b101;
      memory_array[12508] <= 3'b101;
      memory_array[12509] <= 3'b111;
      memory_array[12510] <= 3'b111;
      memory_array[12511] <= 3'b111;
      memory_array[12512] <= 3'b111;
      memory_array[12513] <= 3'b000;
      memory_array[12514] <= 3'b000;
      memory_array[12515] <= 3'b111;
      memory_array[12516] <= 3'b000;
      memory_array[12517] <= 3'b101;
      memory_array[12518] <= 3'b000;
      memory_array[12519] <= 3'b000;
      memory_array[12520] <= 3'b000;
      memory_array[12521] <= 3'b101;
      memory_array[12522] <= 3'b000;
      memory_array[12523] <= 3'b000;
      memory_array[12524] <= 3'b000;
      memory_array[12525] <= 3'b101;
      memory_array[12526] <= 3'b101;
      memory_array[12527] <= 3'b101;
      memory_array[12528] <= 3'b000;
      memory_array[12529] <= 3'b000;
      memory_array[12530] <= 3'b101;
      memory_array[12531] <= 3'b101;
      memory_array[12532] <= 3'b101;
      memory_array[12533] <= 3'b000;
      memory_array[12534] <= 3'b110;
      memory_array[12535] <= 3'b101;
      memory_array[12536] <= 3'b101;
      memory_array[12537] <= 3'b101;
      memory_array[12538] <= 3'b000;
      memory_array[12539] <= 3'b000;
      memory_array[12540] <= 3'b101;
      memory_array[12541] <= 3'b101;
      memory_array[12542] <= 3'b101;
      memory_array[12543] <= 3'b000;
      memory_array[12544] <= 3'b000;
      memory_array[12545] <= 3'b101;
      memory_array[12546] <= 3'b101;
      memory_array[12547] <= 3'b101;
      memory_array[12548] <= 3'b000;
      memory_array[12549] <= 3'b000;
      memory_array[12550] <= 3'b101;
      memory_array[12551] <= 3'b101;
      memory_array[12552] <= 3'b101;
      memory_array[12553] <= 3'b000;
      memory_array[12554] <= 3'b000;
      memory_array[12555] <= 3'b101;
      memory_array[12556] <= 3'b101;
      memory_array[12557] <= 3'b000;
      memory_array[12558] <= 3'b101;
      memory_array[12559] <= 3'b111;
      memory_array[12560] <= 3'b111;
      memory_array[12561] <= 3'b111;
      memory_array[12562] <= 3'b101;
      memory_array[12563] <= 3'b000;
      memory_array[12564] <= 3'b000;
      memory_array[12565] <= 3'b000;
      memory_array[12566] <= 3'b000;
      memory_array[12567] <= 3'b000;
      memory_array[12568] <= 3'b000;
      memory_array[12569] <= 3'b000;
      memory_array[12570] <= 3'b110;
      memory_array[12571] <= 3'b000;
      memory_array[12572] <= 3'b101;
      memory_array[12573] <= 3'b000;
      memory_array[12574] <= 3'b101;
      memory_array[12575] <= 3'b000;
      memory_array[12576] <= 3'b110;
      memory_array[12577] <= 3'b101;
      memory_array[12578] <= 3'b000;
      memory_array[12579] <= 3'b000;
      memory_array[12580] <= 3'b000;
      memory_array[12581] <= 3'b000;
      memory_array[12582] <= 3'b000;
      memory_array[12583] <= 3'b000;
      memory_array[12584] <= 3'b101;
      memory_array[12585] <= 3'b000;
      memory_array[12586] <= 3'b000;
      memory_array[12587] <= 3'b000;
      memory_array[12588] <= 3'b000;
      memory_array[12589] <= 3'b000;
      memory_array[12590] <= 3'b000;
      memory_array[12591] <= 3'b101;
      memory_array[12592] <= 3'b101;
      memory_array[12593] <= 3'b101;
      memory_array[12594] <= 3'b000;
      memory_array[12595] <= 3'b101;
      memory_array[12596] <= 3'b101;
      memory_array[12597] <= 3'b110;
      memory_array[12598] <= 3'b101;
      memory_array[12599] <= 3'b101;
      memory_array[12600] <= 3'b101;
      memory_array[12601] <= 3'b101;
      memory_array[12602] <= 3'b101;
      memory_array[12603] <= 3'b111;
      memory_array[12604] <= 3'b111;
      memory_array[12605] <= 3'b101;
      memory_array[12606] <= 3'b101;
      memory_array[12607] <= 3'b101;
      memory_array[12608] <= 3'b101;
      memory_array[12609] <= 3'b000;
      memory_array[12610] <= 3'b000;
      memory_array[12611] <= 3'b101;
      memory_array[12612] <= 3'b000;
      memory_array[12613] <= 3'b101;
      memory_array[12614] <= 3'b101;
      memory_array[12615] <= 3'b000;
      memory_array[12616] <= 3'b101;
      memory_array[12617] <= 3'b000;
      memory_array[12618] <= 3'b110;
      memory_array[12619] <= 3'b110;
      memory_array[12620] <= 3'b000;
      memory_array[12621] <= 3'b000;
      memory_array[12622] <= 3'b000;
      memory_array[12623] <= 3'b000;
      memory_array[12624] <= 3'b000;
      memory_array[12625] <= 3'b000;
      memory_array[12626] <= 3'b000;
      memory_array[12627] <= 3'b101;
      memory_array[12628] <= 3'b000;
      memory_array[12629] <= 3'b110;
      memory_array[12630] <= 3'b000;
      memory_array[12631] <= 3'b000;
      memory_array[12632] <= 3'b000;
      memory_array[12633] <= 3'b110;
      memory_array[12634] <= 3'b110;
      memory_array[12635] <= 3'b000;
      memory_array[12636] <= 3'b000;
      memory_array[12637] <= 3'b101;
      memory_array[12638] <= 3'b111;
      memory_array[12639] <= 3'b111;
      memory_array[12640] <= 3'b111;
      memory_array[12641] <= 3'b111;
      memory_array[12642] <= 3'b000;
      memory_array[12643] <= 3'b000;
      memory_array[12644] <= 3'b000;
      memory_array[12645] <= 3'b000;
      memory_array[12646] <= 3'b000;
      memory_array[12647] <= 3'b000;
      memory_array[12648] <= 3'b000;
      memory_array[12649] <= 3'b000;
      memory_array[12650] <= 3'b000;
      memory_array[12651] <= 3'b000;
      memory_array[12652] <= 3'b000;
      memory_array[12653] <= 3'b101;
      memory_array[12654] <= 3'b000;
      memory_array[12655] <= 3'b000;
      memory_array[12656] <= 3'b000;
      memory_array[12657] <= 3'b000;
      memory_array[12658] <= 3'b000;
      memory_array[12659] <= 3'b000;
      memory_array[12660] <= 3'b000;
      memory_array[12661] <= 3'b101;
      memory_array[12662] <= 3'b101;
      memory_array[12663] <= 3'b101;
      memory_array[12664] <= 3'b101;
      memory_array[12665] <= 3'b000;
      memory_array[12666] <= 3'b000;
      memory_array[12667] <= 3'b101;
      memory_array[12668] <= 3'b101;
      memory_array[12669] <= 3'b101;
      memory_array[12670] <= 3'b000;
      memory_array[12671] <= 3'b000;
      memory_array[12672] <= 3'b111;
      memory_array[12673] <= 3'b111;
      memory_array[12674] <= 3'b111;
      memory_array[12675] <= 3'b111;
      memory_array[12676] <= 3'b111;
      memory_array[12677] <= 3'b111;
      memory_array[12678] <= 3'b111;
      memory_array[12679] <= 3'b111;
      memory_array[12680] <= 3'b111;
      memory_array[12681] <= 3'b111;
      memory_array[12682] <= 3'b000;
      memory_array[12683] <= 3'b101;
      memory_array[12684] <= 3'b101;
      memory_array[12685] <= 3'b000;
      memory_array[12686] <= 3'b101;
      memory_array[12687] <= 3'b000;
      memory_array[12688] <= 3'b101;
      memory_array[12689] <= 3'b101;
      memory_array[12690] <= 3'b000;
      memory_array[12691] <= 3'b000;
      memory_array[12692] <= 3'b111;
      memory_array[12693] <= 3'b111;
      memory_array[12694] <= 3'b000;
      memory_array[12695] <= 3'b000;
      memory_array[12696] <= 3'b111;
      memory_array[12697] <= 3'b000;
      memory_array[12698] <= 3'b000;
      memory_array[12699] <= 3'b000;
      memory_array[12700] <= 3'b000;
      memory_array[12701] <= 3'b000;
      memory_array[12702] <= 3'b000;
      memory_array[12703] <= 3'b000;
      memory_array[12704] <= 3'b000;
      memory_array[12705] <= 3'b111;
      memory_array[12706] <= 3'b111;
      memory_array[12707] <= 3'b111;
      memory_array[12708] <= 3'b101;
      memory_array[12709] <= 3'b111;
      memory_array[12710] <= 3'b000;
      memory_array[12711] <= 3'b000;
      memory_array[12712] <= 3'b111;
      memory_array[12713] <= 3'b101;
      memory_array[12714] <= 3'b110;
      memory_array[12715] <= 3'b111;
      memory_array[12716] <= 3'b000;
      memory_array[12717] <= 3'b000;
      memory_array[12718] <= 3'b101;
      memory_array[12719] <= 3'b110;
      memory_array[12720] <= 3'b101;
      memory_array[12721] <= 3'b000;
      memory_array[12722] <= 3'b000;
      memory_array[12723] <= 3'b000;
      memory_array[12724] <= 3'b000;
      memory_array[12725] <= 3'b000;
      memory_array[12726] <= 3'b000;
      memory_array[12727] <= 3'b000;
      memory_array[12728] <= 3'b101;
      memory_array[12729] <= 3'b000;
      memory_array[12730] <= 3'b000;
      memory_array[12731] <= 3'b000;
      memory_array[12732] <= 3'b000;
      memory_array[12733] <= 3'b101;
      memory_array[12734] <= 3'b110;
      memory_array[12735] <= 3'b110;
      memory_array[12736] <= 3'b110;
      memory_array[12737] <= 3'b000;
      memory_array[12738] <= 3'b101;
      memory_array[12739] <= 3'b101;
      memory_array[12740] <= 3'b000;
      memory_array[12741] <= 3'b000;
      memory_array[12742] <= 3'b000;
      memory_array[12743] <= 3'b101;
      memory_array[12744] <= 3'b101;
      memory_array[12745] <= 3'b000;
      memory_array[12746] <= 3'b000;
      memory_array[12747] <= 3'b000;
      memory_array[12748] <= 3'b000;
      memory_array[12749] <= 3'b101;
      memory_array[12750] <= 3'b000;
      memory_array[12751] <= 3'b000;
      memory_array[12752] <= 3'b000;
      memory_array[12753] <= 3'b101;
      memory_array[12754] <= 3'b101;
      memory_array[12755] <= 3'b000;
      memory_array[12756] <= 3'b000;
      memory_array[12757] <= 3'b101;
      memory_array[12758] <= 3'b111;
      memory_array[12759] <= 3'b111;
      memory_array[12760] <= 3'b111;
      memory_array[12761] <= 3'b111;
      memory_array[12762] <= 3'b000;
      memory_array[12763] <= 3'b000;
      memory_array[12764] <= 3'b110;
      memory_array[12765] <= 3'b000;
      memory_array[12766] <= 3'b000;
      memory_array[12767] <= 3'b000;
      memory_array[12768] <= 3'b110;
      memory_array[12769] <= 3'b110;
      memory_array[12770] <= 3'b000;
      memory_array[12771] <= 3'b000;
      memory_array[12772] <= 3'b101;
      memory_array[12773] <= 3'b000;
      memory_array[12774] <= 3'b110;
      memory_array[12775] <= 3'b000;
      memory_array[12776] <= 3'b000;
      memory_array[12777] <= 3'b000;
      memory_array[12778] <= 3'b000;
      memory_array[12779] <= 3'b110;
      memory_array[12780] <= 3'b000;
      memory_array[12781] <= 3'b000;
      memory_array[12782] <= 3'b000;
      memory_array[12783] <= 3'b101;
      memory_array[12784] <= 3'b000;
      memory_array[12785] <= 3'b101;
      memory_array[12786] <= 3'b101;
      memory_array[12787] <= 3'b111;
      memory_array[12788] <= 3'b101;
      memory_array[12789] <= 3'b000;
      memory_array[12790] <= 3'b000;
      memory_array[12791] <= 3'b101;
      memory_array[12792] <= 3'b101;
      memory_array[12793] <= 3'b101;
      memory_array[12794] <= 3'b101;
      memory_array[12795] <= 3'b111;
      memory_array[12796] <= 3'b111;
      memory_array[12797] <= 3'b101;
      memory_array[12798] <= 3'b101;
      memory_array[12799] <= 3'b101;
      memory_array[12800] <= 3'b101;
      memory_array[12801] <= 3'b101;
      memory_array[12802] <= 3'b101;
      memory_array[12803] <= 3'b101;
      memory_array[12804] <= 3'b101;
      memory_array[12805] <= 3'b101;
      memory_array[12806] <= 3'b101;
      memory_array[12807] <= 3'b101;
      memory_array[12808] <= 3'b101;
      memory_array[12809] <= 3'b000;
      memory_array[12810] <= 3'b000;
      memory_array[12811] <= 3'b000;
      memory_array[12812] <= 3'b101;
      memory_array[12813] <= 3'b000;
      memory_array[12814] <= 3'b000;
      memory_array[12815] <= 3'b101;
      memory_array[12816] <= 3'b000;
      memory_array[12817] <= 3'b000;
      memory_array[12818] <= 3'b110;
      memory_array[12819] <= 3'b110;
      memory_array[12820] <= 3'b000;
      memory_array[12821] <= 3'b000;
      memory_array[12822] <= 3'b000;
      memory_array[12823] <= 3'b000;
      memory_array[12824] <= 3'b110;
      memory_array[12825] <= 3'b000;
      memory_array[12826] <= 3'b101;
      memory_array[12827] <= 3'b000;
      memory_array[12828] <= 3'b110;
      memory_array[12829] <= 3'b110;
      memory_array[12830] <= 3'b000;
      memory_array[12831] <= 3'b000;
      memory_array[12832] <= 3'b000;
      memory_array[12833] <= 3'b110;
      memory_array[12834] <= 3'b110;
      memory_array[12835] <= 3'b000;
      memory_array[12836] <= 3'b000;
      memory_array[12837] <= 3'b000;
      memory_array[12838] <= 3'b000;
      memory_array[12839] <= 3'b111;
      memory_array[12840] <= 3'b111;
      memory_array[12841] <= 3'b111;
      memory_array[12842] <= 3'b111;
      memory_array[12843] <= 3'b101;
      memory_array[12844] <= 3'b000;
      memory_array[12845] <= 3'b000;
      memory_array[12846] <= 3'b000;
      memory_array[12847] <= 3'b000;
      memory_array[12848] <= 3'b000;
      memory_array[12849] <= 3'b000;
      memory_array[12850] <= 3'b000;
      memory_array[12851] <= 3'b000;
      memory_array[12852] <= 3'b000;
      memory_array[12853] <= 3'b000;
      memory_array[12854] <= 3'b000;
      memory_array[12855] <= 3'b000;
      memory_array[12856] <= 3'b000;
      memory_array[12857] <= 3'b000;
      memory_array[12858] <= 3'b101;
      memory_array[12859] <= 3'b101;
      memory_array[12860] <= 3'b000;
      memory_array[12861] <= 3'b000;
      memory_array[12862] <= 3'b000;
      memory_array[12863] <= 3'b101;
      memory_array[12864] <= 3'b111;
      memory_array[12865] <= 3'b000;
      memory_array[12866] <= 3'b101;
      memory_array[12867] <= 3'b000;
      memory_array[12868] <= 3'b101;
      memory_array[12869] <= 3'b101;
      memory_array[12870] <= 3'b000;
      memory_array[12871] <= 3'b000;
      memory_array[12872] <= 3'b111;
      memory_array[12873] <= 3'b111;
      memory_array[12874] <= 3'b111;
      memory_array[12875] <= 3'b111;
      memory_array[12876] <= 3'b111;
      memory_array[12877] <= 3'b111;
      memory_array[12878] <= 3'b111;
      memory_array[12879] <= 3'b000;
      memory_array[12880] <= 3'b000;
      memory_array[12881] <= 3'b111;
      memory_array[12882] <= 3'b111;
      memory_array[12883] <= 3'b111;
      memory_array[12884] <= 3'b111;
      memory_array[12885] <= 3'b111;
      memory_array[12886] <= 3'b111;
      memory_array[12887] <= 3'b000;
      memory_array[12888] <= 3'b101;
      memory_array[12889] <= 3'b101;
      memory_array[12890] <= 3'b000;
      memory_array[12891] <= 3'b000;
      memory_array[12892] <= 3'b111;
      memory_array[12893] <= 3'b111;
      memory_array[12894] <= 3'b110;
      memory_array[12895] <= 3'b000;
      memory_array[12896] <= 3'b111;
      memory_array[12897] <= 3'b000;
      memory_array[12898] <= 3'b000;
      memory_array[12899] <= 3'b000;
      memory_array[12900] <= 3'b000;
      memory_array[12901] <= 3'b000;
      memory_array[12902] <= 3'b000;
      memory_array[12903] <= 3'b101;
      memory_array[12904] <= 3'b101;
      memory_array[12905] <= 3'b000;
      memory_array[12906] <= 3'b000;
      memory_array[12907] <= 3'b111;
      memory_array[12908] <= 3'b111;
      memory_array[12909] <= 3'b111;
      memory_array[12910] <= 3'b111;
      memory_array[12911] <= 3'b111;
      memory_array[12912] <= 3'b111;
      memory_array[12913] <= 3'b101;
      memory_array[12914] <= 3'b111;
      memory_array[12915] <= 3'b000;
      memory_array[12916] <= 3'b000;
      memory_array[12917] <= 3'b000;
      memory_array[12918] <= 3'b000;
      memory_array[12919] <= 3'b000;
      memory_array[12920] <= 3'b000;
      memory_array[12921] <= 3'b000;
      memory_array[12922] <= 3'b000;
      memory_array[12923] <= 3'b000;
      memory_array[12924] <= 3'b000;
      memory_array[12925] <= 3'b000;
      memory_array[12926] <= 3'b000;
      memory_array[12927] <= 3'b000;
      memory_array[12928] <= 3'b101;
      memory_array[12929] <= 3'b101;
      memory_array[12930] <= 3'b000;
      memory_array[12931] <= 3'b000;
      memory_array[12932] <= 3'b000;
      memory_array[12933] <= 3'b101;
      memory_array[12934] <= 3'b000;
      memory_array[12935] <= 3'b000;
      memory_array[12936] <= 3'b000;
      memory_array[12937] <= 3'b000;
      memory_array[12938] <= 3'b101;
      memory_array[12939] <= 3'b000;
      memory_array[12940] <= 3'b000;
      memory_array[12941] <= 3'b000;
      memory_array[12942] <= 3'b000;
      memory_array[12943] <= 3'b000;
      memory_array[12944] <= 3'b000;
      memory_array[12945] <= 3'b000;
      memory_array[12946] <= 3'b000;
      memory_array[12947] <= 3'b000;
      memory_array[12948] <= 3'b000;
      memory_array[12949] <= 3'b000;
      memory_array[12950] <= 3'b000;
      memory_array[12951] <= 3'b000;
      memory_array[12952] <= 3'b000;
      memory_array[12953] <= 3'b101;
      memory_array[12954] <= 3'b101;
      memory_array[12955] <= 3'b000;
      memory_array[12956] <= 3'b101;
      memory_array[12957] <= 3'b111;
      memory_array[12958] <= 3'b111;
      memory_array[12959] <= 3'b111;
      memory_array[12960] <= 3'b111;
      memory_array[12961] <= 3'b000;
      memory_array[12962] <= 3'b000;
      memory_array[12963] <= 3'b110;
      memory_array[12964] <= 3'b110;
      memory_array[12965] <= 3'b000;
      memory_array[12966] <= 3'b000;
      memory_array[12967] <= 3'b000;
      memory_array[12968] <= 3'b110;
      memory_array[12969] <= 3'b110;
      memory_array[12970] <= 3'b000;
      memory_array[12971] <= 3'b000;
      memory_array[12972] <= 3'b000;
      memory_array[12973] <= 3'b101;
      memory_array[12974] <= 3'b000;
      memory_array[12975] <= 3'b000;
      memory_array[12976] <= 3'b000;
      memory_array[12977] <= 3'b000;
      memory_array[12978] <= 3'b110;
      memory_array[12979] <= 3'b110;
      memory_array[12980] <= 3'b000;
      memory_array[12981] <= 3'b000;
      memory_array[12982] <= 3'b000;
      memory_array[12983] <= 3'b110;
      memory_array[12984] <= 3'b101;
      memory_array[12985] <= 3'b000;
      memory_array[12986] <= 3'b000;
      memory_array[12987] <= 3'b000;
      memory_array[12988] <= 3'b110;
      memory_array[12989] <= 3'b000;
      memory_array[12990] <= 3'b000;
      memory_array[12991] <= 3'b101;
      memory_array[12992] <= 3'b111;
      memory_array[12993] <= 3'b101;
      memory_array[12994] <= 3'b101;
      memory_array[12995] <= 3'b101;
      memory_array[12996] <= 3'b101;
      memory_array[12997] <= 3'b101;
      memory_array[12998] <= 3'b101;
      memory_array[12999] <= 3'b101;
      memory_array[13000] <= 3'b101;
      memory_array[13001] <= 3'b101;
      memory_array[13002] <= 3'b101;
      memory_array[13003] <= 3'b101;
      memory_array[13004] <= 3'b101;
      memory_array[13005] <= 3'b101;
      memory_array[13006] <= 3'b101;
      memory_array[13007] <= 3'b101;
      memory_array[13008] <= 3'b101;
      memory_array[13009] <= 3'b000;
      memory_array[13010] <= 3'b000;
      memory_array[13011] <= 3'b000;
      memory_array[13012] <= 3'b101;
      memory_array[13013] <= 3'b000;
      memory_array[13014] <= 3'b000;
      memory_array[13015] <= 3'b101;
      memory_array[13016] <= 3'b000;
      memory_array[13017] <= 3'b000;
      memory_array[13018] <= 3'b110;
      memory_array[13019] <= 3'b110;
      memory_array[13020] <= 3'b000;
      memory_array[13021] <= 3'b000;
      memory_array[13022] <= 3'b000;
      memory_array[13023] <= 3'b000;
      memory_array[13024] <= 3'b110;
      memory_array[13025] <= 3'b000;
      memory_array[13026] <= 3'b101;
      memory_array[13027] <= 3'b000;
      memory_array[13028] <= 3'b110;
      memory_array[13029] <= 3'b110;
      memory_array[13030] <= 3'b000;
      memory_array[13031] <= 3'b000;
      memory_array[13032] <= 3'b000;
      memory_array[13033] <= 3'b110;
      memory_array[13034] <= 3'b110;
      memory_array[13035] <= 3'b000;
      memory_array[13036] <= 3'b000;
      memory_array[13037] <= 3'b000;
      memory_array[13038] <= 3'b000;
      memory_array[13039] <= 3'b111;
      memory_array[13040] <= 3'b111;
      memory_array[13041] <= 3'b111;
      memory_array[13042] <= 3'b111;
      memory_array[13043] <= 3'b101;
      memory_array[13044] <= 3'b000;
      memory_array[13045] <= 3'b000;
      memory_array[13046] <= 3'b000;
      memory_array[13047] <= 3'b000;
      memory_array[13048] <= 3'b000;
      memory_array[13049] <= 3'b000;
      memory_array[13050] <= 3'b000;
      memory_array[13051] <= 3'b000;
      memory_array[13052] <= 3'b000;
      memory_array[13053] <= 3'b000;
      memory_array[13054] <= 3'b000;
      memory_array[13055] <= 3'b000;
      memory_array[13056] <= 3'b000;
      memory_array[13057] <= 3'b000;
      memory_array[13058] <= 3'b101;
      memory_array[13059] <= 3'b101;
      memory_array[13060] <= 3'b000;
      memory_array[13061] <= 3'b000;
      memory_array[13062] <= 3'b000;
      memory_array[13063] <= 3'b101;
      memory_array[13064] <= 3'b111;
      memory_array[13065] <= 3'b000;
      memory_array[13066] <= 3'b101;
      memory_array[13067] <= 3'b000;
      memory_array[13068] <= 3'b101;
      memory_array[13069] <= 3'b101;
      memory_array[13070] <= 3'b000;
      memory_array[13071] <= 3'b000;
      memory_array[13072] <= 3'b111;
      memory_array[13073] <= 3'b111;
      memory_array[13074] <= 3'b111;
      memory_array[13075] <= 3'b111;
      memory_array[13076] <= 3'b111;
      memory_array[13077] <= 3'b111;
      memory_array[13078] <= 3'b111;
      memory_array[13079] <= 3'b000;
      memory_array[13080] <= 3'b000;
      memory_array[13081] <= 3'b111;
      memory_array[13082] <= 3'b111;
      memory_array[13083] <= 3'b111;
      memory_array[13084] <= 3'b111;
      memory_array[13085] <= 3'b111;
      memory_array[13086] <= 3'b111;
      memory_array[13087] <= 3'b000;
      memory_array[13088] <= 3'b101;
      memory_array[13089] <= 3'b101;
      memory_array[13090] <= 3'b000;
      memory_array[13091] <= 3'b000;
      memory_array[13092] <= 3'b111;
      memory_array[13093] <= 3'b111;
      memory_array[13094] <= 3'b110;
      memory_array[13095] <= 3'b000;
      memory_array[13096] <= 3'b111;
      memory_array[13097] <= 3'b000;
      memory_array[13098] <= 3'b000;
      memory_array[13099] <= 3'b000;
      memory_array[13100] <= 3'b000;
      memory_array[13101] <= 3'b000;
      memory_array[13102] <= 3'b000;
      memory_array[13103] <= 3'b101;
      memory_array[13104] <= 3'b101;
      memory_array[13105] <= 3'b000;
      memory_array[13106] <= 3'b000;
      memory_array[13107] <= 3'b111;
      memory_array[13108] <= 3'b111;
      memory_array[13109] <= 3'b111;
      memory_array[13110] <= 3'b111;
      memory_array[13111] <= 3'b111;
      memory_array[13112] <= 3'b111;
      memory_array[13113] <= 3'b101;
      memory_array[13114] <= 3'b111;
      memory_array[13115] <= 3'b000;
      memory_array[13116] <= 3'b000;
      memory_array[13117] <= 3'b000;
      memory_array[13118] <= 3'b000;
      memory_array[13119] <= 3'b000;
      memory_array[13120] <= 3'b000;
      memory_array[13121] <= 3'b000;
      memory_array[13122] <= 3'b000;
      memory_array[13123] <= 3'b000;
      memory_array[13124] <= 3'b000;
      memory_array[13125] <= 3'b000;
      memory_array[13126] <= 3'b000;
      memory_array[13127] <= 3'b000;
      memory_array[13128] <= 3'b101;
      memory_array[13129] <= 3'b101;
      memory_array[13130] <= 3'b000;
      memory_array[13131] <= 3'b000;
      memory_array[13132] <= 3'b000;
      memory_array[13133] <= 3'b101;
      memory_array[13134] <= 3'b000;
      memory_array[13135] <= 3'b000;
      memory_array[13136] <= 3'b000;
      memory_array[13137] <= 3'b000;
      memory_array[13138] <= 3'b101;
      memory_array[13139] <= 3'b000;
      memory_array[13140] <= 3'b000;
      memory_array[13141] <= 3'b000;
      memory_array[13142] <= 3'b000;
      memory_array[13143] <= 3'b000;
      memory_array[13144] <= 3'b000;
      memory_array[13145] <= 3'b000;
      memory_array[13146] <= 3'b000;
      memory_array[13147] <= 3'b000;
      memory_array[13148] <= 3'b000;
      memory_array[13149] <= 3'b000;
      memory_array[13150] <= 3'b000;
      memory_array[13151] <= 3'b000;
      memory_array[13152] <= 3'b000;
      memory_array[13153] <= 3'b101;
      memory_array[13154] <= 3'b101;
      memory_array[13155] <= 3'b000;
      memory_array[13156] <= 3'b101;
      memory_array[13157] <= 3'b111;
      memory_array[13158] <= 3'b111;
      memory_array[13159] <= 3'b111;
      memory_array[13160] <= 3'b111;
      memory_array[13161] <= 3'b000;
      memory_array[13162] <= 3'b000;
      memory_array[13163] <= 3'b110;
      memory_array[13164] <= 3'b110;
      memory_array[13165] <= 3'b000;
      memory_array[13166] <= 3'b000;
      memory_array[13167] <= 3'b000;
      memory_array[13168] <= 3'b110;
      memory_array[13169] <= 3'b110;
      memory_array[13170] <= 3'b000;
      memory_array[13171] <= 3'b000;
      memory_array[13172] <= 3'b000;
      memory_array[13173] <= 3'b101;
      memory_array[13174] <= 3'b000;
      memory_array[13175] <= 3'b000;
      memory_array[13176] <= 3'b000;
      memory_array[13177] <= 3'b000;
      memory_array[13178] <= 3'b110;
      memory_array[13179] <= 3'b110;
      memory_array[13180] <= 3'b000;
      memory_array[13181] <= 3'b000;
      memory_array[13182] <= 3'b000;
      memory_array[13183] <= 3'b110;
      memory_array[13184] <= 3'b101;
      memory_array[13185] <= 3'b000;
      memory_array[13186] <= 3'b000;
      memory_array[13187] <= 3'b000;
      memory_array[13188] <= 3'b110;
      memory_array[13189] <= 3'b000;
      memory_array[13190] <= 3'b000;
      memory_array[13191] <= 3'b101;
      memory_array[13192] <= 3'b111;
      memory_array[13193] <= 3'b101;
      memory_array[13194] <= 3'b101;
      memory_array[13195] <= 3'b101;
      memory_array[13196] <= 3'b101;
      memory_array[13197] <= 3'b101;
      memory_array[13198] <= 3'b101;
      memory_array[13199] <= 3'b101;
      memory_array[13200] <= 3'b101;
      memory_array[13201] <= 3'b101;
      memory_array[13202] <= 3'b101;
      memory_array[13203] <= 3'b111;
      memory_array[13204] <= 3'b111;
      memory_array[13205] <= 3'b101;
      memory_array[13206] <= 3'b101;
      memory_array[13207] <= 3'b101;
      memory_array[13208] <= 3'b101;
      memory_array[13209] <= 3'b000;
      memory_array[13210] <= 3'b000;
      memory_array[13211] <= 3'b000;
      memory_array[13212] <= 3'b000;
      memory_array[13213] <= 3'b000;
      memory_array[13214] <= 3'b000;
      memory_array[13215] <= 3'b000;
      memory_array[13216] <= 3'b000;
      memory_array[13217] <= 3'b000;
      memory_array[13218] <= 3'b000;
      memory_array[13219] <= 3'b000;
      memory_array[13220] <= 3'b000;
      memory_array[13221] <= 3'b000;
      memory_array[13222] <= 3'b000;
      memory_array[13223] <= 3'b000;
      memory_array[13224] <= 3'b000;
      memory_array[13225] <= 3'b000;
      memory_array[13226] <= 3'b000;
      memory_array[13227] <= 3'b000;
      memory_array[13228] <= 3'b000;
      memory_array[13229] <= 3'b000;
      memory_array[13230] <= 3'b000;
      memory_array[13231] <= 3'b000;
      memory_array[13232] <= 3'b000;
      memory_array[13233] <= 3'b000;
      memory_array[13234] <= 3'b000;
      memory_array[13235] <= 3'b000;
      memory_array[13236] <= 3'b000;
      memory_array[13237] <= 3'b000;
      memory_array[13238] <= 3'b000;
      memory_array[13239] <= 3'b000;
      memory_array[13240] <= 3'b101;
      memory_array[13241] <= 3'b111;
      memory_array[13242] <= 3'b111;
      memory_array[13243] <= 3'b111;
      memory_array[13244] <= 3'b111;
      memory_array[13245] <= 3'b101;
      memory_array[13246] <= 3'b000;
      memory_array[13247] <= 3'b000;
      memory_array[13248] <= 3'b000;
      memory_array[13249] <= 3'b000;
      memory_array[13250] <= 3'b000;
      memory_array[13251] <= 3'b000;
      memory_array[13252] <= 3'b000;
      memory_array[13253] <= 3'b000;
      memory_array[13254] <= 3'b000;
      memory_array[13255] <= 3'b000;
      memory_array[13256] <= 3'b000;
      memory_array[13257] <= 3'b000;
      memory_array[13258] <= 3'b101;
      memory_array[13259] <= 3'b000;
      memory_array[13260] <= 3'b000;
      memory_array[13261] <= 3'b000;
      memory_array[13262] <= 3'b000;
      memory_array[13263] <= 3'b000;
      memory_array[13264] <= 3'b000;
      memory_array[13265] <= 3'b000;
      memory_array[13266] <= 3'b000;
      memory_array[13267] <= 3'b000;
      memory_array[13268] <= 3'b000;
      memory_array[13269] <= 3'b000;
      memory_array[13270] <= 3'b000;
      memory_array[13271] <= 3'b000;
      memory_array[13272] <= 3'b000;
      memory_array[13273] <= 3'b000;
      memory_array[13274] <= 3'b000;
      memory_array[13275] <= 3'b000;
      memory_array[13276] <= 3'b000;
      memory_array[13277] <= 3'b000;
      memory_array[13278] <= 3'b000;
      memory_array[13279] <= 3'b000;
      memory_array[13280] <= 3'b000;
      memory_array[13281] <= 3'b111;
      memory_array[13282] <= 3'b111;
      memory_array[13283] <= 3'b111;
      memory_array[13284] <= 3'b000;
      memory_array[13285] <= 3'b000;
      memory_array[13286] <= 3'b000;
      memory_array[13287] <= 3'b111;
      memory_array[13288] <= 3'b111;
      memory_array[13289] <= 3'b000;
      memory_array[13290] <= 3'b000;
      memory_array[13291] <= 3'b000;
      memory_array[13292] <= 3'b111;
      memory_array[13293] <= 3'b111;
      memory_array[13294] <= 3'b111;
      memory_array[13295] <= 3'b111;
      memory_array[13296] <= 3'b000;
      memory_array[13297] <= 3'b000;
      memory_array[13298] <= 3'b101;
      memory_array[13299] <= 3'b101;
      memory_array[13300] <= 3'b000;
      memory_array[13301] <= 3'b000;
      memory_array[13302] <= 3'b000;
      memory_array[13303] <= 3'b000;
      memory_array[13304] <= 3'b000;
      memory_array[13305] <= 3'b000;
      memory_array[13306] <= 3'b000;
      memory_array[13307] <= 3'b000;
      memory_array[13308] <= 3'b101;
      memory_array[13309] <= 3'b101;
      memory_array[13310] <= 3'b111;
      memory_array[13311] <= 3'b111;
      memory_array[13312] <= 3'b111;
      memory_array[13313] <= 3'b111;
      memory_array[13314] <= 3'b101;
      memory_array[13315] <= 3'b000;
      memory_array[13316] <= 3'b111;
      memory_array[13317] <= 3'b000;
      memory_array[13318] <= 3'b101;
      memory_array[13319] <= 3'b101;
      memory_array[13320] <= 3'b000;
      memory_array[13321] <= 3'b000;
      memory_array[13322] <= 3'b000;
      memory_array[13323] <= 3'b000;
      memory_array[13324] <= 3'b101;
      memory_array[13325] <= 3'b000;
      memory_array[13326] <= 3'b000;
      memory_array[13327] <= 3'b000;
      memory_array[13328] <= 3'b101;
      memory_array[13329] <= 3'b000;
      memory_array[13330] <= 3'b000;
      memory_array[13331] <= 3'b000;
      memory_array[13332] <= 3'b000;
      memory_array[13333] <= 3'b101;
      memory_array[13334] <= 3'b101;
      memory_array[13335] <= 3'b000;
      memory_array[13336] <= 3'b000;
      memory_array[13337] <= 3'b000;
      memory_array[13338] <= 3'b110;
      memory_array[13339] <= 3'b000;
      memory_array[13340] <= 3'b000;
      memory_array[13341] <= 3'b000;
      memory_array[13342] <= 3'b000;
      memory_array[13343] <= 3'b000;
      memory_array[13344] <= 3'b000;
      memory_array[13345] <= 3'b000;
      memory_array[13346] <= 3'b000;
      memory_array[13347] <= 3'b000;
      memory_array[13348] <= 3'b000;
      memory_array[13349] <= 3'b000;
      memory_array[13350] <= 3'b000;
      memory_array[13351] <= 3'b000;
      memory_array[13352] <= 3'b000;
      memory_array[13353] <= 3'b000;
      memory_array[13354] <= 3'b101;
      memory_array[13355] <= 3'b111;
      memory_array[13356] <= 3'b111;
      memory_array[13357] <= 3'b111;
      memory_array[13358] <= 3'b111;
      memory_array[13359] <= 3'b101;
      memory_array[13360] <= 3'b000;
      memory_array[13361] <= 3'b000;
      memory_array[13362] <= 3'b000;
      memory_array[13363] <= 3'b000;
      memory_array[13364] <= 3'b000;
      memory_array[13365] <= 3'b000;
      memory_array[13366] <= 3'b000;
      memory_array[13367] <= 3'b000;
      memory_array[13368] <= 3'b000;
      memory_array[13369] <= 3'b000;
      memory_array[13370] <= 3'b000;
      memory_array[13371] <= 3'b000;
      memory_array[13372] <= 3'b000;
      memory_array[13373] <= 3'b000;
      memory_array[13374] <= 3'b000;
      memory_array[13375] <= 3'b000;
      memory_array[13376] <= 3'b000;
      memory_array[13377] <= 3'b000;
      memory_array[13378] <= 3'b000;
      memory_array[13379] <= 3'b000;
      memory_array[13380] <= 3'b000;
      memory_array[13381] <= 3'b000;
      memory_array[13382] <= 3'b000;
      memory_array[13383] <= 3'b000;
      memory_array[13384] <= 3'b000;
      memory_array[13385] <= 3'b000;
      memory_array[13386] <= 3'b000;
      memory_array[13387] <= 3'b000;
      memory_array[13388] <= 3'b000;
      memory_array[13389] <= 3'b000;
      memory_array[13390] <= 3'b000;
      memory_array[13391] <= 3'b101;
      memory_array[13392] <= 3'b101;
      memory_array[13393] <= 3'b101;
      memory_array[13394] <= 3'b101;
      memory_array[13395] <= 3'b111;
      memory_array[13396] <= 3'b111;
      memory_array[13397] <= 3'b101;
      memory_array[13398] <= 3'b101;
      memory_array[13399] <= 3'b101;
      memory_array[13400] <= 3'b101;
      memory_array[13401] <= 3'b000;
      memory_array[13402] <= 3'b000;
      memory_array[13403] <= 3'b110;
      memory_array[13404] <= 3'b110;
      memory_array[13405] <= 3'b000;
      memory_array[13406] <= 3'b000;
      memory_array[13407] <= 3'b101;
      memory_array[13408] <= 3'b101;
      memory_array[13409] <= 3'b000;
      memory_array[13410] <= 3'b000;
      memory_array[13411] <= 3'b101;
      memory_array[13412] <= 3'b101;
      memory_array[13413] <= 3'b101;
      memory_array[13414] <= 3'b111;
      memory_array[13415] <= 3'b111;
      memory_array[13416] <= 3'b111;
      memory_array[13417] <= 3'b111;
      memory_array[13418] <= 3'b111;
      memory_array[13419] <= 3'b101;
      memory_array[13420] <= 3'b101;
      memory_array[13421] <= 3'b101;
      memory_array[13422] <= 3'b101;
      memory_array[13423] <= 3'b101;
      memory_array[13424] <= 3'b111;
      memory_array[13425] <= 3'b111;
      memory_array[13426] <= 3'b111;
      memory_array[13427] <= 3'b111;
      memory_array[13428] <= 3'b111;
      memory_array[13429] <= 3'b101;
      memory_array[13430] <= 3'b101;
      memory_array[13431] <= 3'b101;
      memory_array[13432] <= 3'b101;
      memory_array[13433] <= 3'b101;
      memory_array[13434] <= 3'b111;
      memory_array[13435] <= 3'b111;
      memory_array[13436] <= 3'b111;
      memory_array[13437] <= 3'b111;
      memory_array[13438] <= 3'b111;
      memory_array[13439] <= 3'b101;
      memory_array[13440] <= 3'b101;
      memory_array[13441] <= 3'b101;
      memory_array[13442] <= 3'b111;
      memory_array[13443] <= 3'b111;
      memory_array[13444] <= 3'b111;
      memory_array[13445] <= 3'b111;
      memory_array[13446] <= 3'b111;
      memory_array[13447] <= 3'b000;
      memory_array[13448] <= 3'b000;
      memory_array[13449] <= 3'b000;
      memory_array[13450] <= 3'b000;
      memory_array[13451] <= 3'b000;
      memory_array[13452] <= 3'b000;
      memory_array[13453] <= 3'b101;
      memory_array[13454] <= 3'b000;
      memory_array[13455] <= 3'b000;
      memory_array[13456] <= 3'b000;
      memory_array[13457] <= 3'b000;
      memory_array[13458] <= 3'b000;
      memory_array[13459] <= 3'b101;
      memory_array[13460] <= 3'b000;
      memory_array[13461] <= 3'b000;
      memory_array[13462] <= 3'b000;
      memory_array[13463] <= 3'b101;
      memory_array[13464] <= 3'b101;
      memory_array[13465] <= 3'b101;
      memory_array[13466] <= 3'b101;
      memory_array[13467] <= 3'b101;
      memory_array[13468] <= 3'b111;
      memory_array[13469] <= 3'b111;
      memory_array[13470] <= 3'b111;
      memory_array[13471] <= 3'b111;
      memory_array[13472] <= 3'b101;
      memory_array[13473] <= 3'b111;
      memory_array[13474] <= 3'b101;
      memory_array[13475] <= 3'b101;
      memory_array[13476] <= 3'b000;
      memory_array[13477] <= 3'b000;
      memory_array[13478] <= 3'b000;
      memory_array[13479] <= 3'b000;
      memory_array[13480] <= 3'b000;
      memory_array[13481] <= 3'b000;
      memory_array[13482] <= 3'b000;
      memory_array[13483] <= 3'b101;
      memory_array[13484] <= 3'b000;
      memory_array[13485] <= 3'b000;
      memory_array[13486] <= 3'b000;
      memory_array[13487] <= 3'b111;
      memory_array[13488] <= 3'b111;
      memory_array[13489] <= 3'b000;
      memory_array[13490] <= 3'b000;
      memory_array[13491] <= 3'b000;
      memory_array[13492] <= 3'b000;
      memory_array[13493] <= 3'b101;
      memory_array[13494] <= 3'b101;
      memory_array[13495] <= 3'b111;
      memory_array[13496] <= 3'b101;
      memory_array[13497] <= 3'b000;
      memory_array[13498] <= 3'b110;
      memory_array[13499] <= 3'b110;
      memory_array[13500] <= 3'b000;
      memory_array[13501] <= 3'b000;
      memory_array[13502] <= 3'b000;
      memory_array[13503] <= 3'b110;
      memory_array[13504] <= 3'b101;
      memory_array[13505] <= 3'b000;
      memory_array[13506] <= 3'b000;
      memory_array[13507] <= 3'b000;
      memory_array[13508] <= 3'b110;
      memory_array[13509] <= 3'b110;
      memory_array[13510] <= 3'b000;
      memory_array[13511] <= 3'b000;
      memory_array[13512] <= 3'b000;
      memory_array[13513] <= 3'b101;
      memory_array[13514] <= 3'b000;
      memory_array[13515] <= 3'b000;
      memory_array[13516] <= 3'b000;
      memory_array[13517] <= 3'b000;
      memory_array[13518] <= 3'b000;
      memory_array[13519] <= 3'b000;
      memory_array[13520] <= 3'b000;
      memory_array[13521] <= 3'b000;
      memory_array[13522] <= 3'b000;
      memory_array[13523] <= 3'b000;
      memory_array[13524] <= 3'b000;
      memory_array[13525] <= 3'b000;
      memory_array[13526] <= 3'b000;
      memory_array[13527] <= 3'b000;
      memory_array[13528] <= 3'b000;
      memory_array[13529] <= 3'b000;
      memory_array[13530] <= 3'b000;
      memory_array[13531] <= 3'b000;
      memory_array[13532] <= 3'b000;
      memory_array[13533] <= 3'b000;
      memory_array[13534] <= 3'b000;
      memory_array[13535] <= 3'b000;
      memory_array[13536] <= 3'b000;
      memory_array[13537] <= 3'b000;
      memory_array[13538] <= 3'b000;
      memory_array[13539] <= 3'b000;
      memory_array[13540] <= 3'b000;
      memory_array[13541] <= 3'b000;
      memory_array[13542] <= 3'b000;
      memory_array[13543] <= 3'b110;
      memory_array[13544] <= 3'b000;
      memory_array[13545] <= 3'b000;
      memory_array[13546] <= 3'b000;
      memory_array[13547] <= 3'b000;
      memory_array[13548] <= 3'b000;
      memory_array[13549] <= 3'b000;
      memory_array[13550] <= 3'b000;
      memory_array[13551] <= 3'b000;
      memory_array[13552] <= 3'b101;
      memory_array[13553] <= 3'b111;
      memory_array[13554] <= 3'b111;
      memory_array[13555] <= 3'b111;
      memory_array[13556] <= 3'b111;
      memory_array[13557] <= 3'b111;
      memory_array[13558] <= 3'b101;
      memory_array[13559] <= 3'b101;
      memory_array[13560] <= 3'b101;
      memory_array[13561] <= 3'b111;
      memory_array[13562] <= 3'b111;
      memory_array[13563] <= 3'b111;
      memory_array[13564] <= 3'b111;
      memory_array[13565] <= 3'b111;
      memory_array[13566] <= 3'b101;
      memory_array[13567] <= 3'b101;
      memory_array[13568] <= 3'b101;
      memory_array[13569] <= 3'b101;
      memory_array[13570] <= 3'b101;
      memory_array[13571] <= 3'b111;
      memory_array[13572] <= 3'b111;
      memory_array[13573] <= 3'b111;
      memory_array[13574] <= 3'b111;
      memory_array[13575] <= 3'b111;
      memory_array[13576] <= 3'b101;
      memory_array[13577] <= 3'b101;
      memory_array[13578] <= 3'b101;
      memory_array[13579] <= 3'b101;
      memory_array[13580] <= 3'b101;
      memory_array[13581] <= 3'b111;
      memory_array[13582] <= 3'b111;
      memory_array[13583] <= 3'b111;
      memory_array[13584] <= 3'b111;
      memory_array[13585] <= 3'b111;
      memory_array[13586] <= 3'b101;
      memory_array[13587] <= 3'b101;
      memory_array[13588] <= 3'b101;
      memory_array[13589] <= 3'b000;
      memory_array[13590] <= 3'b000;
      memory_array[13591] <= 3'b101;
      memory_array[13592] <= 3'b101;
      memory_array[13593] <= 3'b110;
      memory_array[13594] <= 3'b110;
      memory_array[13595] <= 3'b000;
      memory_array[13596] <= 3'b000;
      memory_array[13597] <= 3'b000;
      memory_array[13598] <= 3'b110;
      memory_array[13599] <= 3'b101;
      memory_array[13600] <= 3'b101;
      memory_array[13601] <= 3'b110;
      memory_array[13602] <= 3'b110;
      memory_array[13603] <= 3'b000;
      memory_array[13604] <= 3'b000;
      memory_array[13605] <= 3'b110;
      memory_array[13606] <= 3'b110;
      memory_array[13607] <= 3'b101;
      memory_array[13608] <= 3'b101;
      memory_array[13609] <= 3'b000;
      memory_array[13610] <= 3'b000;
      memory_array[13611] <= 3'b101;
      memory_array[13612] <= 3'b101;
      memory_array[13613] <= 3'b101;
      memory_array[13614] <= 3'b111;
      memory_array[13615] <= 3'b111;
      memory_array[13616] <= 3'b111;
      memory_array[13617] <= 3'b111;
      memory_array[13618] <= 3'b111;
      memory_array[13619] <= 3'b101;
      memory_array[13620] <= 3'b101;
      memory_array[13621] <= 3'b101;
      memory_array[13622] <= 3'b101;
      memory_array[13623] <= 3'b101;
      memory_array[13624] <= 3'b111;
      memory_array[13625] <= 3'b111;
      memory_array[13626] <= 3'b111;
      memory_array[13627] <= 3'b111;
      memory_array[13628] <= 3'b111;
      memory_array[13629] <= 3'b101;
      memory_array[13630] <= 3'b101;
      memory_array[13631] <= 3'b101;
      memory_array[13632] <= 3'b101;
      memory_array[13633] <= 3'b101;
      memory_array[13634] <= 3'b111;
      memory_array[13635] <= 3'b111;
      memory_array[13636] <= 3'b111;
      memory_array[13637] <= 3'b111;
      memory_array[13638] <= 3'b111;
      memory_array[13639] <= 3'b101;
      memory_array[13640] <= 3'b101;
      memory_array[13641] <= 3'b000;
      memory_array[13642] <= 3'b111;
      memory_array[13643] <= 3'b111;
      memory_array[13644] <= 3'b111;
      memory_array[13645] <= 3'b111;
      memory_array[13646] <= 3'b111;
      memory_array[13647] <= 3'b111;
      memory_array[13648] <= 3'b101;
      memory_array[13649] <= 3'b000;
      memory_array[13650] <= 3'b000;
      memory_array[13651] <= 3'b000;
      memory_array[13652] <= 3'b101;
      memory_array[13653] <= 3'b000;
      memory_array[13654] <= 3'b000;
      memory_array[13655] <= 3'b000;
      memory_array[13656] <= 3'b000;
      memory_array[13657] <= 3'b000;
      memory_array[13658] <= 3'b000;
      memory_array[13659] <= 3'b000;
      memory_array[13660] <= 3'b000;
      memory_array[13661] <= 3'b101;
      memory_array[13662] <= 3'b000;
      memory_array[13663] <= 3'b000;
      memory_array[13664] <= 3'b000;
      memory_array[13665] <= 3'b000;
      memory_array[13666] <= 3'b000;
      memory_array[13667] <= 3'b000;
      memory_array[13668] <= 3'b000;
      memory_array[13669] <= 3'b000;
      memory_array[13670] <= 3'b101;
      memory_array[13671] <= 3'b101;
      memory_array[13672] <= 3'b101;
      memory_array[13673] <= 3'b000;
      memory_array[13674] <= 3'b101;
      memory_array[13675] <= 3'b101;
      memory_array[13676] <= 3'b101;
      memory_array[13677] <= 3'b000;
      memory_array[13678] <= 3'b000;
      memory_array[13679] <= 3'b000;
      memory_array[13680] <= 3'b101;
      memory_array[13681] <= 3'b000;
      memory_array[13682] <= 3'b101;
      memory_array[13683] <= 3'b000;
      memory_array[13684] <= 3'b000;
      memory_array[13685] <= 3'b000;
      memory_array[13686] <= 3'b000;
      memory_array[13687] <= 3'b000;
      memory_array[13688] <= 3'b000;
      memory_array[13689] <= 3'b000;
      memory_array[13690] <= 3'b000;
      memory_array[13691] <= 3'b101;
      memory_array[13692] <= 3'b111;
      memory_array[13693] <= 3'b111;
      memory_array[13694] <= 3'b101;
      memory_array[13695] <= 3'b110;
      memory_array[13696] <= 3'b110;
      memory_array[13697] <= 3'b110;
      memory_array[13698] <= 3'b000;
      memory_array[13699] <= 3'b000;
      memory_array[13700] <= 3'b110;
      memory_array[13701] <= 3'b110;
      memory_array[13702] <= 3'b110;
      memory_array[13703] <= 3'b000;
      memory_array[13704] <= 3'b000;
      memory_array[13705] <= 3'b000;
      memory_array[13706] <= 3'b000;
      memory_array[13707] <= 3'b000;
      memory_array[13708] <= 3'b000;
      memory_array[13709] <= 3'b000;
      memory_array[13710] <= 3'b101;
      memory_array[13711] <= 3'b101;
      memory_array[13712] <= 3'b101;
      memory_array[13713] <= 3'b101;
      memory_array[13714] <= 3'b101;
      memory_array[13715] <= 3'b101;
      memory_array[13716] <= 3'b101;
      memory_array[13717] <= 3'b101;
      memory_array[13718] <= 3'b000;
      memory_array[13719] <= 3'b000;
      memory_array[13720] <= 3'b101;
      memory_array[13721] <= 3'b101;
      memory_array[13722] <= 3'b101;
      memory_array[13723] <= 3'b000;
      memory_array[13724] <= 3'b000;
      memory_array[13725] <= 3'b000;
      memory_array[13726] <= 3'b101;
      memory_array[13727] <= 3'b101;
      memory_array[13728] <= 3'b101;
      memory_array[13729] <= 3'b101;
      memory_array[13730] <= 3'b101;
      memory_array[13731] <= 3'b101;
      memory_array[13732] <= 3'b110;
      memory_array[13733] <= 3'b111;
      memory_array[13734] <= 3'b110;
      memory_array[13735] <= 3'b110;
      memory_array[13736] <= 3'b000;
      memory_array[13737] <= 3'b000;
      memory_array[13738] <= 3'b000;
      memory_array[13739] <= 3'b000;
      memory_array[13740] <= 3'b000;
      memory_array[13741] <= 3'b110;
      memory_array[13742] <= 3'b110;
      memory_array[13743] <= 3'b000;
      memory_array[13744] <= 3'b000;
      memory_array[13745] <= 3'b000;
      memory_array[13746] <= 3'b000;
      memory_array[13747] <= 3'b000;
      memory_array[13748] <= 3'b000;
      memory_array[13749] <= 3'b000;
      memory_array[13750] <= 3'b000;
      memory_array[13751] <= 3'b101;
      memory_array[13752] <= 3'b111;
      memory_array[13753] <= 3'b111;
      memory_array[13754] <= 3'b111;
      memory_array[13755] <= 3'b111;
      memory_array[13756] <= 3'b111;
      memory_array[13757] <= 3'b101;
      memory_array[13758] <= 3'b000;
      memory_array[13759] <= 3'b101;
      memory_array[13760] <= 3'b101;
      memory_array[13761] <= 3'b111;
      memory_array[13762] <= 3'b111;
      memory_array[13763] <= 3'b111;
      memory_array[13764] <= 3'b111;
      memory_array[13765] <= 3'b111;
      memory_array[13766] <= 3'b101;
      memory_array[13767] <= 3'b101;
      memory_array[13768] <= 3'b101;
      memory_array[13769] <= 3'b101;
      memory_array[13770] <= 3'b101;
      memory_array[13771] <= 3'b111;
      memory_array[13772] <= 3'b111;
      memory_array[13773] <= 3'b111;
      memory_array[13774] <= 3'b111;
      memory_array[13775] <= 3'b111;
      memory_array[13776] <= 3'b101;
      memory_array[13777] <= 3'b101;
      memory_array[13778] <= 3'b101;
      memory_array[13779] <= 3'b101;
      memory_array[13780] <= 3'b101;
      memory_array[13781] <= 3'b111;
      memory_array[13782] <= 3'b111;
      memory_array[13783] <= 3'b111;
      memory_array[13784] <= 3'b111;
      memory_array[13785] <= 3'b111;
      memory_array[13786] <= 3'b101;
      memory_array[13787] <= 3'b101;
      memory_array[13788] <= 3'b101;
      memory_array[13789] <= 3'b000;
      memory_array[13790] <= 3'b000;
      memory_array[13791] <= 3'b101;
      memory_array[13792] <= 3'b110;
      memory_array[13793] <= 3'b000;
      memory_array[13794] <= 3'b000;
      memory_array[13795] <= 3'b110;
      memory_array[13796] <= 3'b110;
      memory_array[13797] <= 3'b110;
      memory_array[13798] <= 3'b000;
      memory_array[13799] <= 3'b101;
      memory_array[13800] <= 3'b000;
      memory_array[13801] <= 3'b000;
      memory_array[13802] <= 3'b000;
      memory_array[13803] <= 3'b110;
      memory_array[13804] <= 3'b110;
      memory_array[13805] <= 3'b000;
      memory_array[13806] <= 3'b000;
      memory_array[13807] <= 3'b000;
      memory_array[13808] <= 3'b101;
      memory_array[13809] <= 3'b000;
      memory_array[13810] <= 3'b000;
      memory_array[13811] <= 3'b101;
      memory_array[13812] <= 3'b101;
      memory_array[13813] <= 3'b101;
      memory_array[13814] <= 3'b111;
      memory_array[13815] <= 3'b111;
      memory_array[13816] <= 3'b111;
      memory_array[13817] <= 3'b111;
      memory_array[13818] <= 3'b111;
      memory_array[13819] <= 3'b101;
      memory_array[13820] <= 3'b101;
      memory_array[13821] <= 3'b101;
      memory_array[13822] <= 3'b101;
      memory_array[13823] <= 3'b101;
      memory_array[13824] <= 3'b111;
      memory_array[13825] <= 3'b111;
      memory_array[13826] <= 3'b111;
      memory_array[13827] <= 3'b111;
      memory_array[13828] <= 3'b111;
      memory_array[13829] <= 3'b101;
      memory_array[13830] <= 3'b101;
      memory_array[13831] <= 3'b101;
      memory_array[13832] <= 3'b101;
      memory_array[13833] <= 3'b101;
      memory_array[13834] <= 3'b111;
      memory_array[13835] <= 3'b111;
      memory_array[13836] <= 3'b111;
      memory_array[13837] <= 3'b111;
      memory_array[13838] <= 3'b111;
      memory_array[13839] <= 3'b101;
      memory_array[13840] <= 3'b101;
      memory_array[13841] <= 3'b101;
      memory_array[13842] <= 3'b101;
      memory_array[13843] <= 3'b111;
      memory_array[13844] <= 3'b111;
      memory_array[13845] <= 3'b111;
      memory_array[13846] <= 3'b111;
      memory_array[13847] <= 3'b111;
      memory_array[13848] <= 3'b111;
      memory_array[13849] <= 3'b000;
      memory_array[13850] <= 3'b000;
      memory_array[13851] <= 3'b000;
      memory_array[13852] <= 3'b000;
      memory_array[13853] <= 3'b101;
      memory_array[13854] <= 3'b000;
      memory_array[13855] <= 3'b000;
      memory_array[13856] <= 3'b000;
      memory_array[13857] <= 3'b000;
      memory_array[13858] <= 3'b000;
      memory_array[13859] <= 3'b000;
      memory_array[13860] <= 3'b000;
      memory_array[13861] <= 3'b000;
      memory_array[13862] <= 3'b000;
      memory_array[13863] <= 3'b000;
      memory_array[13864] <= 3'b000;
      memory_array[13865] <= 3'b000;
      memory_array[13866] <= 3'b000;
      memory_array[13867] <= 3'b000;
      memory_array[13868] <= 3'b000;
      memory_array[13869] <= 3'b000;
      memory_array[13870] <= 3'b000;
      memory_array[13871] <= 3'b000;
      memory_array[13872] <= 3'b101;
      memory_array[13873] <= 3'b000;
      memory_array[13874] <= 3'b101;
      memory_array[13875] <= 3'b000;
      memory_array[13876] <= 3'b000;
      memory_array[13877] <= 3'b000;
      memory_array[13878] <= 3'b000;
      memory_array[13879] <= 3'b101;
      memory_array[13880] <= 3'b000;
      memory_array[13881] <= 3'b000;
      memory_array[13882] <= 3'b000;
      memory_array[13883] <= 3'b101;
      memory_array[13884] <= 3'b000;
      memory_array[13885] <= 3'b000;
      memory_array[13886] <= 3'b000;
      memory_array[13887] <= 3'b000;
      memory_array[13888] <= 3'b000;
      memory_array[13889] <= 3'b000;
      memory_array[13890] <= 3'b101;
      memory_array[13891] <= 3'b000;
      memory_array[13892] <= 3'b000;
      memory_array[13893] <= 3'b000;
      memory_array[13894] <= 3'b101;
      memory_array[13895] <= 3'b000;
      memory_array[13896] <= 3'b000;
      memory_array[13897] <= 3'b000;
      memory_array[13898] <= 3'b110;
      memory_array[13899] <= 3'b110;
      memory_array[13900] <= 3'b000;
      memory_array[13901] <= 3'b000;
      memory_array[13902] <= 3'b000;
      memory_array[13903] <= 3'b000;
      memory_array[13904] <= 3'b101;
      memory_array[13905] <= 3'b000;
      memory_array[13906] <= 3'b000;
      memory_array[13907] <= 3'b101;
      memory_array[13908] <= 3'b101;
      memory_array[13909] <= 3'b101;
      memory_array[13910] <= 3'b000;
      memory_array[13911] <= 3'b000;
      memory_array[13912] <= 3'b000;
      memory_array[13913] <= 3'b101;
      memory_array[13914] <= 3'b101;
      memory_array[13915] <= 3'b000;
      memory_array[13916] <= 3'b000;
      memory_array[13917] <= 3'b000;
      memory_array[13918] <= 3'b101;
      memory_array[13919] <= 3'b101;
      memory_array[13920] <= 3'b000;
      memory_array[13921] <= 3'b000;
      memory_array[13922] <= 3'b000;
      memory_array[13923] <= 3'b101;
      memory_array[13924] <= 3'b101;
      memory_array[13925] <= 3'b101;
      memory_array[13926] <= 3'b111;
      memory_array[13927] <= 3'b110;
      memory_array[13928] <= 3'b110;
      memory_array[13929] <= 3'b110;
      memory_array[13930] <= 3'b111;
      memory_array[13931] <= 3'b111;
      memory_array[13932] <= 3'b111;
      memory_array[13933] <= 3'b101;
      memory_array[13934] <= 3'b101;
      memory_array[13935] <= 3'b000;
      memory_array[13936] <= 3'b000;
      memory_array[13937] <= 3'b000;
      memory_array[13938] <= 3'b000;
      memory_array[13939] <= 3'b110;
      memory_array[13940] <= 3'b000;
      memory_array[13941] <= 3'b000;
      memory_array[13942] <= 3'b000;
      memory_array[13943] <= 3'b000;
      memory_array[13944] <= 3'b000;
      memory_array[13945] <= 3'b000;
      memory_array[13946] <= 3'b000;
      memory_array[13947] <= 3'b000;
      memory_array[13948] <= 3'b000;
      memory_array[13949] <= 3'b000;
      memory_array[13950] <= 3'b101;
      memory_array[13951] <= 3'b111;
      memory_array[13952] <= 3'b111;
      memory_array[13953] <= 3'b111;
      memory_array[13954] <= 3'b111;
      memory_array[13955] <= 3'b111;
      memory_array[13956] <= 3'b111;
      memory_array[13957] <= 3'b000;
      memory_array[13958] <= 3'b101;
      memory_array[13959] <= 3'b101;
      memory_array[13960] <= 3'b101;
      memory_array[13961] <= 3'b111;
      memory_array[13962] <= 3'b111;
      memory_array[13963] <= 3'b111;
      memory_array[13964] <= 3'b111;
      memory_array[13965] <= 3'b111;
      memory_array[13966] <= 3'b101;
      memory_array[13967] <= 3'b101;
      memory_array[13968] <= 3'b101;
      memory_array[13969] <= 3'b101;
      memory_array[13970] <= 3'b101;
      memory_array[13971] <= 3'b111;
      memory_array[13972] <= 3'b111;
      memory_array[13973] <= 3'b111;
      memory_array[13974] <= 3'b111;
      memory_array[13975] <= 3'b111;
      memory_array[13976] <= 3'b101;
      memory_array[13977] <= 3'b101;
      memory_array[13978] <= 3'b101;
      memory_array[13979] <= 3'b101;
      memory_array[13980] <= 3'b101;
      memory_array[13981] <= 3'b111;
      memory_array[13982] <= 3'b111;
      memory_array[13983] <= 3'b111;
      memory_array[13984] <= 3'b111;
      memory_array[13985] <= 3'b111;
      memory_array[13986] <= 3'b101;
      memory_array[13987] <= 3'b101;
      memory_array[13988] <= 3'b101;
      memory_array[13989] <= 3'b000;
      memory_array[13990] <= 3'b000;
      memory_array[13991] <= 3'b101;
      memory_array[13992] <= 3'b000;
      memory_array[13993] <= 3'b110;
      memory_array[13994] <= 3'b110;
      memory_array[13995] <= 3'b000;
      memory_array[13996] <= 3'b000;
      memory_array[13997] <= 3'b000;
      memory_array[13998] <= 3'b110;
      memory_array[13999] <= 3'b110;
      memory_array[14000] <= 3'b101;
      memory_array[14001] <= 3'b101;
      memory_array[14002] <= 3'b101;
      memory_array[14003] <= 3'b101;
      memory_array[14004] <= 3'b101;
      memory_array[14005] <= 3'b101;
      memory_array[14006] <= 3'b101;
      memory_array[14007] <= 3'b101;
      memory_array[14008] <= 3'b101;
      memory_array[14009] <= 3'b000;
      memory_array[14010] <= 3'b000;
      memory_array[14011] <= 3'b101;
      memory_array[14012] <= 3'b101;
      memory_array[14013] <= 3'b101;
      memory_array[14014] <= 3'b111;
      memory_array[14015] <= 3'b111;
      memory_array[14016] <= 3'b111;
      memory_array[14017] <= 3'b111;
      memory_array[14018] <= 3'b111;
      memory_array[14019] <= 3'b101;
      memory_array[14020] <= 3'b101;
      memory_array[14021] <= 3'b101;
      memory_array[14022] <= 3'b101;
      memory_array[14023] <= 3'b101;
      memory_array[14024] <= 3'b111;
      memory_array[14025] <= 3'b111;
      memory_array[14026] <= 3'b111;
      memory_array[14027] <= 3'b111;
      memory_array[14028] <= 3'b111;
      memory_array[14029] <= 3'b101;
      memory_array[14030] <= 3'b101;
      memory_array[14031] <= 3'b101;
      memory_array[14032] <= 3'b101;
      memory_array[14033] <= 3'b101;
      memory_array[14034] <= 3'b111;
      memory_array[14035] <= 3'b111;
      memory_array[14036] <= 3'b111;
      memory_array[14037] <= 3'b111;
      memory_array[14038] <= 3'b111;
      memory_array[14039] <= 3'b101;
      memory_array[14040] <= 3'b101;
      memory_array[14041] <= 3'b101;
      memory_array[14042] <= 3'b000;
      memory_array[14043] <= 3'b101;
      memory_array[14044] <= 3'b111;
      memory_array[14045] <= 3'b111;
      memory_array[14046] <= 3'b111;
      memory_array[14047] <= 3'b111;
      memory_array[14048] <= 3'b111;
      memory_array[14049] <= 3'b101;
      memory_array[14050] <= 3'b000;
      memory_array[14051] <= 3'b000;
      memory_array[14052] <= 3'b101;
      memory_array[14053] <= 3'b000;
      memory_array[14054] <= 3'b000;
      memory_array[14055] <= 3'b000;
      memory_array[14056] <= 3'b000;
      memory_array[14057] <= 3'b000;
      memory_array[14058] <= 3'b000;
      memory_array[14059] <= 3'b000;
      memory_array[14060] <= 3'b000;
      memory_array[14061] <= 3'b101;
      memory_array[14062] <= 3'b000;
      memory_array[14063] <= 3'b000;
      memory_array[14064] <= 3'b000;
      memory_array[14065] <= 3'b000;
      memory_array[14066] <= 3'b000;
      memory_array[14067] <= 3'b000;
      memory_array[14068] <= 3'b000;
      memory_array[14069] <= 3'b000;
      memory_array[14070] <= 3'b000;
      memory_array[14071] <= 3'b000;
      memory_array[14072] <= 3'b101;
      memory_array[14073] <= 3'b101;
      memory_array[14074] <= 3'b101;
      memory_array[14075] <= 3'b101;
      memory_array[14076] <= 3'b101;
      memory_array[14077] <= 3'b101;
      memory_array[14078] <= 3'b000;
      memory_array[14079] <= 3'b000;
      memory_array[14080] <= 3'b101;
      memory_array[14081] <= 3'b101;
      memory_array[14082] <= 3'b101;
      memory_array[14083] <= 3'b000;
      memory_array[14084] <= 3'b000;
      memory_array[14085] <= 3'b000;
      memory_array[14086] <= 3'b000;
      memory_array[14087] <= 3'b000;
      memory_array[14088] <= 3'b000;
      memory_array[14089] <= 3'b000;
      memory_array[14090] <= 3'b000;
      memory_array[14091] <= 3'b000;
      memory_array[14092] <= 3'b000;
      memory_array[14093] <= 3'b000;
      memory_array[14094] <= 3'b000;
      memory_array[14095] <= 3'b000;
      memory_array[14096] <= 3'b000;
      memory_array[14097] <= 3'b000;
      memory_array[14098] <= 3'b000;
      memory_array[14099] <= 3'b000;
      memory_array[14100] <= 3'b101;
      memory_array[14101] <= 3'b101;
      memory_array[14102] <= 3'b101;
      memory_array[14103] <= 3'b000;
      memory_array[14104] <= 3'b000;
      memory_array[14105] <= 3'b101;
      memory_array[14106] <= 3'b101;
      memory_array[14107] <= 3'b101;
      memory_array[14108] <= 3'b000;
      memory_array[14109] <= 3'b000;
      memory_array[14110] <= 3'b000;
      memory_array[14111] <= 3'b000;
      memory_array[14112] <= 3'b000;
      memory_array[14113] <= 3'b000;
      memory_array[14114] <= 3'b000;
      memory_array[14115] <= 3'b000;
      memory_array[14116] <= 3'b000;
      memory_array[14117] <= 3'b000;
      memory_array[14118] <= 3'b000;
      memory_array[14119] <= 3'b000;
      memory_array[14120] <= 3'b000;
      memory_array[14121] <= 3'b000;
      memory_array[14122] <= 3'b000;
      memory_array[14123] <= 3'b000;
      memory_array[14124] <= 3'b000;
      memory_array[14125] <= 3'b000;
      memory_array[14126] <= 3'b000;
      memory_array[14127] <= 3'b101;
      memory_array[14128] <= 3'b101;
      memory_array[14129] <= 3'b101;
      memory_array[14130] <= 3'b101;
      memory_array[14131] <= 3'b101;
      memory_array[14132] <= 3'b101;
      memory_array[14133] <= 3'b101;
      memory_array[14134] <= 3'b000;
      memory_array[14135] <= 3'b000;
      memory_array[14136] <= 3'b000;
      memory_array[14137] <= 3'b000;
      memory_array[14138] <= 3'b000;
      memory_array[14139] <= 3'b000;
      memory_array[14140] <= 3'b110;
      memory_array[14141] <= 3'b000;
      memory_array[14142] <= 3'b000;
      memory_array[14143] <= 3'b000;
      memory_array[14144] <= 3'b000;
      memory_array[14145] <= 3'b000;
      memory_array[14146] <= 3'b000;
      memory_array[14147] <= 3'b110;
      memory_array[14148] <= 3'b000;
      memory_array[14149] <= 3'b000;
      memory_array[14150] <= 3'b111;
      memory_array[14151] <= 3'b111;
      memory_array[14152] <= 3'b111;
      memory_array[14153] <= 3'b111;
      memory_array[14154] <= 3'b111;
      memory_array[14155] <= 3'b111;
      memory_array[14156] <= 3'b101;
      memory_array[14157] <= 3'b101;
      memory_array[14158] <= 3'b101;
      memory_array[14159] <= 3'b101;
      memory_array[14160] <= 3'b101;
      memory_array[14161] <= 3'b111;
      memory_array[14162] <= 3'b111;
      memory_array[14163] <= 3'b111;
      memory_array[14164] <= 3'b111;
      memory_array[14165] <= 3'b111;
      memory_array[14166] <= 3'b101;
      memory_array[14167] <= 3'b101;
      memory_array[14168] <= 3'b101;
      memory_array[14169] <= 3'b101;
      memory_array[14170] <= 3'b101;
      memory_array[14171] <= 3'b111;
      memory_array[14172] <= 3'b111;
      memory_array[14173] <= 3'b111;
      memory_array[14174] <= 3'b111;
      memory_array[14175] <= 3'b111;
      memory_array[14176] <= 3'b101;
      memory_array[14177] <= 3'b101;
      memory_array[14178] <= 3'b101;
      memory_array[14179] <= 3'b101;
      memory_array[14180] <= 3'b101;
      memory_array[14181] <= 3'b111;
      memory_array[14182] <= 3'b111;
      memory_array[14183] <= 3'b111;
      memory_array[14184] <= 3'b111;
      memory_array[14185] <= 3'b111;
      memory_array[14186] <= 3'b101;
      memory_array[14187] <= 3'b101;
      memory_array[14188] <= 3'b101;
      memory_array[14189] <= 3'b000;
      memory_array[14190] <= 3'b000;
      memory_array[14191] <= 3'b101;
      memory_array[14192] <= 3'b101;
      memory_array[14193] <= 3'b101;
      memory_array[14194] <= 3'b101;
      memory_array[14195] <= 3'b101;
      memory_array[14196] <= 3'b101;
      memory_array[14197] <= 3'b101;
      memory_array[14198] <= 3'b101;
      memory_array[14199] <= 3'b101;
      memory_array[14200] <= 3'b101;
      memory_array[14201] <= 3'b101;
      memory_array[14202] <= 3'b101;
      memory_array[14203] <= 3'b101;
      memory_array[14204] <= 3'b101;
      memory_array[14205] <= 3'b101;
      memory_array[14206] <= 3'b101;
      memory_array[14207] <= 3'b101;
      memory_array[14208] <= 3'b101;
      memory_array[14209] <= 3'b000;
      memory_array[14210] <= 3'b000;
      memory_array[14211] <= 3'b101;
      memory_array[14212] <= 3'b101;
      memory_array[14213] <= 3'b101;
      memory_array[14214] <= 3'b111;
      memory_array[14215] <= 3'b111;
      memory_array[14216] <= 3'b111;
      memory_array[14217] <= 3'b111;
      memory_array[14218] <= 3'b111;
      memory_array[14219] <= 3'b101;
      memory_array[14220] <= 3'b101;
      memory_array[14221] <= 3'b101;
      memory_array[14222] <= 3'b101;
      memory_array[14223] <= 3'b101;
      memory_array[14224] <= 3'b111;
      memory_array[14225] <= 3'b111;
      memory_array[14226] <= 3'b111;
      memory_array[14227] <= 3'b111;
      memory_array[14228] <= 3'b111;
      memory_array[14229] <= 3'b101;
      memory_array[14230] <= 3'b101;
      memory_array[14231] <= 3'b101;
      memory_array[14232] <= 3'b101;
      memory_array[14233] <= 3'b101;
      memory_array[14234] <= 3'b111;
      memory_array[14235] <= 3'b111;
      memory_array[14236] <= 3'b111;
      memory_array[14237] <= 3'b111;
      memory_array[14238] <= 3'b111;
      memory_array[14239] <= 3'b101;
      memory_array[14240] <= 3'b101;
      memory_array[14241] <= 3'b101;
      memory_array[14242] <= 3'b101;
      memory_array[14243] <= 3'b101;
      memory_array[14244] <= 3'b111;
      memory_array[14245] <= 3'b111;
      memory_array[14246] <= 3'b111;
      memory_array[14247] <= 3'b111;
      memory_array[14248] <= 3'b111;
      memory_array[14249] <= 3'b101;
      memory_array[14250] <= 3'b000;
      memory_array[14251] <= 3'b000;
      memory_array[14252] <= 3'b000;
      memory_array[14253] <= 3'b000;
      memory_array[14254] <= 3'b000;
      memory_array[14255] <= 3'b000;
      memory_array[14256] <= 3'b000;
      memory_array[14257] <= 3'b000;
      memory_array[14258] <= 3'b000;
      memory_array[14259] <= 3'b000;
      memory_array[14260] <= 3'b000;
      memory_array[14261] <= 3'b101;
      memory_array[14262] <= 3'b000;
      memory_array[14263] <= 3'b000;
      memory_array[14264] <= 3'b000;
      memory_array[14265] <= 3'b000;
      memory_array[14266] <= 3'b000;
      memory_array[14267] <= 3'b000;
      memory_array[14268] <= 3'b000;
      memory_array[14269] <= 3'b000;
      memory_array[14270] <= 3'b000;
      memory_array[14271] <= 3'b000;
      memory_array[14272] <= 3'b000;
      memory_array[14273] <= 3'b000;
      memory_array[14274] <= 3'b000;
      memory_array[14275] <= 3'b000;
      memory_array[14276] <= 3'b101;
      memory_array[14277] <= 3'b101;
      memory_array[14278] <= 3'b000;
      memory_array[14279] <= 3'b000;
      memory_array[14280] <= 3'b000;
      memory_array[14281] <= 3'b000;
      memory_array[14282] <= 3'b101;
      memory_array[14283] <= 3'b111;
      memory_array[14284] <= 3'b111;
      memory_array[14285] <= 3'b111;
      memory_array[14286] <= 3'b101;
      memory_array[14287] <= 3'b101;
      memory_array[14288] <= 3'b101;
      memory_array[14289] <= 3'b101;
      memory_array[14290] <= 3'b101;
      memory_array[14291] <= 3'b101;
      memory_array[14292] <= 3'b101;
      memory_array[14293] <= 3'b101;
      memory_array[14294] <= 3'b000;
      memory_array[14295] <= 3'b000;
      memory_array[14296] <= 3'b101;
      memory_array[14297] <= 3'b101;
      memory_array[14298] <= 3'b000;
      memory_array[14299] <= 3'b000;
      memory_array[14300] <= 3'b000;
      memory_array[14301] <= 3'b000;
      memory_array[14302] <= 3'b000;
      memory_array[14303] <= 3'b000;
      memory_array[14304] <= 3'b000;
      memory_array[14305] <= 3'b101;
      memory_array[14306] <= 3'b000;
      memory_array[14307] <= 3'b101;
      memory_array[14308] <= 3'b111;
      memory_array[14309] <= 3'b101;
      memory_array[14310] <= 3'b101;
      memory_array[14311] <= 3'b101;
      memory_array[14312] <= 3'b101;
      memory_array[14313] <= 3'b000;
      memory_array[14314] <= 3'b000;
      memory_array[14315] <= 3'b101;
      memory_array[14316] <= 3'b101;
      memory_array[14317] <= 3'b101;
      memory_array[14318] <= 3'b000;
      memory_array[14319] <= 3'b000;
      memory_array[14320] <= 3'b000;
      memory_array[14321] <= 3'b000;
      memory_array[14322] <= 3'b101;
      memory_array[14323] <= 3'b000;
      memory_array[14324] <= 3'b000;
      memory_array[14325] <= 3'b101;
      memory_array[14326] <= 3'b101;
      memory_array[14327] <= 3'b101;
      memory_array[14328] <= 3'b000;
      memory_array[14329] <= 3'b000;
      memory_array[14330] <= 3'b000;
      memory_array[14331] <= 3'b000;
      memory_array[14332] <= 3'b000;
      memory_array[14333] <= 3'b000;
      memory_array[14334] <= 3'b000;
      memory_array[14335] <= 3'b110;
      memory_array[14336] <= 3'b110;
      memory_array[14337] <= 3'b110;
      memory_array[14338] <= 3'b000;
      memory_array[14339] <= 3'b000;
      memory_array[14340] <= 3'b000;
      memory_array[14341] <= 3'b000;
      memory_array[14342] <= 3'b000;
      memory_array[14343] <= 3'b000;
      memory_array[14344] <= 3'b000;
      memory_array[14345] <= 3'b000;
      memory_array[14346] <= 3'b110;
      memory_array[14347] <= 3'b101;
      memory_array[14348] <= 3'b000;
      memory_array[14349] <= 3'b000;
      memory_array[14350] <= 3'b111;
      memory_array[14351] <= 3'b111;
      memory_array[14352] <= 3'b111;
      memory_array[14353] <= 3'b111;
      memory_array[14354] <= 3'b111;
      memory_array[14355] <= 3'b101;
      memory_array[14356] <= 3'b101;
      memory_array[14357] <= 3'b101;
      memory_array[14358] <= 3'b101;
      memory_array[14359] <= 3'b101;
      memory_array[14360] <= 3'b101;
      memory_array[14361] <= 3'b111;
      memory_array[14362] <= 3'b111;
      memory_array[14363] <= 3'b111;
      memory_array[14364] <= 3'b111;
      memory_array[14365] <= 3'b111;
      memory_array[14366] <= 3'b101;
      memory_array[14367] <= 3'b101;
      memory_array[14368] <= 3'b101;
      memory_array[14369] <= 3'b101;
      memory_array[14370] <= 3'b101;
      memory_array[14371] <= 3'b111;
      memory_array[14372] <= 3'b111;
      memory_array[14373] <= 3'b111;
      memory_array[14374] <= 3'b111;
      memory_array[14375] <= 3'b111;
      memory_array[14376] <= 3'b101;
      memory_array[14377] <= 3'b101;
      memory_array[14378] <= 3'b101;
      memory_array[14379] <= 3'b101;
      memory_array[14380] <= 3'b101;
      memory_array[14381] <= 3'b111;
      memory_array[14382] <= 3'b111;
      memory_array[14383] <= 3'b111;
      memory_array[14384] <= 3'b111;
      memory_array[14385] <= 3'b111;
      memory_array[14386] <= 3'b101;
      memory_array[14387] <= 3'b101;
      memory_array[14388] <= 3'b101;
      memory_array[14389] <= 3'b000;
      memory_array[14390] <= 3'b000;
      memory_array[14391] <= 3'b101;
      memory_array[14392] <= 3'b101;
      memory_array[14393] <= 3'b101;
      memory_array[14394] <= 3'b101;
      memory_array[14395] <= 3'b101;
      memory_array[14396] <= 3'b101;
      memory_array[14397] <= 3'b101;
      memory_array[14398] <= 3'b101;
      memory_array[14399] <= 3'b101;
      memory_array[14400] <= 3'b000;
      memory_array[14401] <= 3'b000;
      memory_array[14402] <= 3'b000;
      memory_array[14403] <= 3'b110;
      memory_array[14404] <= 3'b110;
      memory_array[14405] <= 3'b000;
      memory_array[14406] <= 3'b000;
      memory_array[14407] <= 3'b000;
      memory_array[14408] <= 3'b101;
      memory_array[14409] <= 3'b000;
      memory_array[14410] <= 3'b000;
      memory_array[14411] <= 3'b101;
      memory_array[14412] <= 3'b101;
      memory_array[14413] <= 3'b101;
      memory_array[14414] <= 3'b111;
      memory_array[14415] <= 3'b111;
      memory_array[14416] <= 3'b111;
      memory_array[14417] <= 3'b111;
      memory_array[14418] <= 3'b111;
      memory_array[14419] <= 3'b101;
      memory_array[14420] <= 3'b101;
      memory_array[14421] <= 3'b101;
      memory_array[14422] <= 3'b101;
      memory_array[14423] <= 3'b101;
      memory_array[14424] <= 3'b111;
      memory_array[14425] <= 3'b111;
      memory_array[14426] <= 3'b111;
      memory_array[14427] <= 3'b111;
      memory_array[14428] <= 3'b111;
      memory_array[14429] <= 3'b101;
      memory_array[14430] <= 3'b101;
      memory_array[14431] <= 3'b101;
      memory_array[14432] <= 3'b101;
      memory_array[14433] <= 3'b101;
      memory_array[14434] <= 3'b111;
      memory_array[14435] <= 3'b111;
      memory_array[14436] <= 3'b111;
      memory_array[14437] <= 3'b111;
      memory_array[14438] <= 3'b111;
      memory_array[14439] <= 3'b101;
      memory_array[14440] <= 3'b101;
      memory_array[14441] <= 3'b101;
      memory_array[14442] <= 3'b101;
      memory_array[14443] <= 3'b101;
      memory_array[14444] <= 3'b111;
      memory_array[14445] <= 3'b111;
      memory_array[14446] <= 3'b111;
      memory_array[14447] <= 3'b111;
      memory_array[14448] <= 3'b111;
      memory_array[14449] <= 3'b101;
      memory_array[14450] <= 3'b000;
      memory_array[14451] <= 3'b000;
      memory_array[14452] <= 3'b000;
      memory_array[14453] <= 3'b000;
      memory_array[14454] <= 3'b101;
      memory_array[14455] <= 3'b000;
      memory_array[14456] <= 3'b000;
      memory_array[14457] <= 3'b000;
      memory_array[14458] <= 3'b000;
      memory_array[14459] <= 3'b000;
      memory_array[14460] <= 3'b000;
      memory_array[14461] <= 3'b000;
      memory_array[14462] <= 3'b000;
      memory_array[14463] <= 3'b000;
      memory_array[14464] <= 3'b000;
      memory_array[14465] <= 3'b000;
      memory_array[14466] <= 3'b000;
      memory_array[14467] <= 3'b000;
      memory_array[14468] <= 3'b000;
      memory_array[14469] <= 3'b000;
      memory_array[14470] <= 3'b000;
      memory_array[14471] <= 3'b000;
      memory_array[14472] <= 3'b000;
      memory_array[14473] <= 3'b000;
      memory_array[14474] <= 3'b000;
      memory_array[14475] <= 3'b000;
      memory_array[14476] <= 3'b000;
      memory_array[14477] <= 3'b000;
      memory_array[14478] <= 3'b000;
      memory_array[14479] <= 3'b000;
      memory_array[14480] <= 3'b000;
      memory_array[14481] <= 3'b111;
      memory_array[14482] <= 3'b111;
      memory_array[14483] <= 3'b101;
      memory_array[14484] <= 3'b101;
      memory_array[14485] <= 3'b101;
      memory_array[14486] <= 3'b101;
      memory_array[14487] <= 3'b101;
      memory_array[14488] <= 3'b101;
      memory_array[14489] <= 3'b101;
      memory_array[14490] <= 3'b000;
      memory_array[14491] <= 3'b000;
      memory_array[14492] <= 3'b000;
      memory_array[14493] <= 3'b101;
      memory_array[14494] <= 3'b101;
      memory_array[14495] <= 3'b000;
      memory_array[14496] <= 3'b000;
      memory_array[14497] <= 3'b000;
      memory_array[14498] <= 3'b000;
      memory_array[14499] <= 3'b000;
      memory_array[14500] <= 3'b000;
      memory_array[14501] <= 3'b101;
      memory_array[14502] <= 3'b111;
      memory_array[14503] <= 3'b111;
      memory_array[14504] <= 3'b111;
      memory_array[14505] <= 3'b101;
      memory_array[14506] <= 3'b101;
      memory_array[14507] <= 3'b101;
      memory_array[14508] <= 3'b101;
      memory_array[14509] <= 3'b101;
      memory_array[14510] <= 3'b000;
      memory_array[14511] <= 3'b000;
      memory_array[14512] <= 3'b101;
      memory_array[14513] <= 3'b101;
      memory_array[14514] <= 3'b101;
      memory_array[14515] <= 3'b101;
      memory_array[14516] <= 3'b000;
      memory_array[14517] <= 3'b000;
      memory_array[14518] <= 3'b000;
      memory_array[14519] <= 3'b101;
      memory_array[14520] <= 3'b000;
      memory_array[14521] <= 3'b000;
      memory_array[14522] <= 3'b101;
      memory_array[14523] <= 3'b101;
      memory_array[14524] <= 3'b101;
      memory_array[14525] <= 3'b101;
      memory_array[14526] <= 3'b101;
      memory_array[14527] <= 3'b101;
      memory_array[14528] <= 3'b101;
      memory_array[14529] <= 3'b101;
      memory_array[14530] <= 3'b101;
      memory_array[14531] <= 3'b000;
      memory_array[14532] <= 3'b000;
      memory_array[14533] <= 3'b000;
      memory_array[14534] <= 3'b110;
      memory_array[14535] <= 3'b000;
      memory_array[14536] <= 3'b000;
      memory_array[14537] <= 3'b000;
      memory_array[14538] <= 3'b000;
      memory_array[14539] <= 3'b000;
      memory_array[14540] <= 3'b000;
      memory_array[14541] <= 3'b000;
      memory_array[14542] <= 3'b000;
      memory_array[14543] <= 3'b000;
      memory_array[14544] <= 3'b000;
      memory_array[14545] <= 3'b000;
      memory_array[14546] <= 3'b000;
      memory_array[14547] <= 3'b000;
      memory_array[14548] <= 3'b101;
      memory_array[14549] <= 3'b000;
      memory_array[14550] <= 3'b111;
      memory_array[14551] <= 3'b111;
      memory_array[14552] <= 3'b111;
      memory_array[14553] <= 3'b111;
      memory_array[14554] <= 3'b111;
      memory_array[14555] <= 3'b101;
      memory_array[14556] <= 3'b101;
      memory_array[14557] <= 3'b101;
      memory_array[14558] <= 3'b101;
      memory_array[14559] <= 3'b101;
      memory_array[14560] <= 3'b101;
      memory_array[14561] <= 3'b111;
      memory_array[14562] <= 3'b111;
      memory_array[14563] <= 3'b111;
      memory_array[14564] <= 3'b111;
      memory_array[14565] <= 3'b111;
      memory_array[14566] <= 3'b101;
      memory_array[14567] <= 3'b101;
      memory_array[14568] <= 3'b101;
      memory_array[14569] <= 3'b101;
      memory_array[14570] <= 3'b101;
      memory_array[14571] <= 3'b111;
      memory_array[14572] <= 3'b111;
      memory_array[14573] <= 3'b111;
      memory_array[14574] <= 3'b111;
      memory_array[14575] <= 3'b111;
      memory_array[14576] <= 3'b101;
      memory_array[14577] <= 3'b101;
      memory_array[14578] <= 3'b101;
      memory_array[14579] <= 3'b101;
      memory_array[14580] <= 3'b101;
      memory_array[14581] <= 3'b111;
      memory_array[14582] <= 3'b111;
      memory_array[14583] <= 3'b111;
      memory_array[14584] <= 3'b111;
      memory_array[14585] <= 3'b111;
      memory_array[14586] <= 3'b101;
      memory_array[14587] <= 3'b101;
      memory_array[14588] <= 3'b101;
      memory_array[14589] <= 3'b000;
      memory_array[14590] <= 3'b000;
      memory_array[14591] <= 3'b101;
      memory_array[14592] <= 3'b000;
      memory_array[14593] <= 3'b110;
      memory_array[14594] <= 3'b110;
      memory_array[14595] <= 3'b000;
      memory_array[14596] <= 3'b000;
      memory_array[14597] <= 3'b000;
      memory_array[14598] <= 3'b110;
      memory_array[14599] <= 3'b110;
      memory_array[14600] <= 3'b101;
      memory_array[14601] <= 3'b110;
      memory_array[14602] <= 3'b110;
      memory_array[14603] <= 3'b000;
      memory_array[14604] <= 3'b000;
      memory_array[14605] <= 3'b110;
      memory_array[14606] <= 3'b110;
      memory_array[14607] <= 3'b101;
      memory_array[14608] <= 3'b101;
      memory_array[14609] <= 3'b000;
      memory_array[14610] <= 3'b000;
      memory_array[14611] <= 3'b101;
      memory_array[14612] <= 3'b101;
      memory_array[14613] <= 3'b101;
      memory_array[14614] <= 3'b111;
      memory_array[14615] <= 3'b111;
      memory_array[14616] <= 3'b111;
      memory_array[14617] <= 3'b111;
      memory_array[14618] <= 3'b111;
      memory_array[14619] <= 3'b101;
      memory_array[14620] <= 3'b101;
      memory_array[14621] <= 3'b101;
      memory_array[14622] <= 3'b101;
      memory_array[14623] <= 3'b101;
      memory_array[14624] <= 3'b111;
      memory_array[14625] <= 3'b111;
      memory_array[14626] <= 3'b111;
      memory_array[14627] <= 3'b111;
      memory_array[14628] <= 3'b111;
      memory_array[14629] <= 3'b101;
      memory_array[14630] <= 3'b101;
      memory_array[14631] <= 3'b101;
      memory_array[14632] <= 3'b101;
      memory_array[14633] <= 3'b101;
      memory_array[14634] <= 3'b111;
      memory_array[14635] <= 3'b111;
      memory_array[14636] <= 3'b111;
      memory_array[14637] <= 3'b111;
      memory_array[14638] <= 3'b111;
      memory_array[14639] <= 3'b101;
      memory_array[14640] <= 3'b101;
      memory_array[14641] <= 3'b101;
      memory_array[14642] <= 3'b101;
      memory_array[14643] <= 3'b101;
      memory_array[14644] <= 3'b111;
      memory_array[14645] <= 3'b111;
      memory_array[14646] <= 3'b111;
      memory_array[14647] <= 3'b111;
      memory_array[14648] <= 3'b111;
      memory_array[14649] <= 3'b101;
      memory_array[14650] <= 3'b000;
      memory_array[14651] <= 3'b000;
      memory_array[14652] <= 3'b000;
      memory_array[14653] <= 3'b000;
      memory_array[14654] <= 3'b000;
      memory_array[14655] <= 3'b101;
      memory_array[14656] <= 3'b000;
      memory_array[14657] <= 3'b000;
      memory_array[14658] <= 3'b000;
      memory_array[14659] <= 3'b000;
      memory_array[14660] <= 3'b000;
      memory_array[14661] <= 3'b000;
      memory_array[14662] <= 3'b000;
      memory_array[14663] <= 3'b000;
      memory_array[14664] <= 3'b000;
      memory_array[14665] <= 3'b000;
      memory_array[14666] <= 3'b000;
      memory_array[14667] <= 3'b110;
      memory_array[14668] <= 3'b000;
      memory_array[14669] <= 3'b000;
      memory_array[14670] <= 3'b000;
      memory_array[14671] <= 3'b000;
      memory_array[14672] <= 3'b000;
      memory_array[14673] <= 3'b000;
      memory_array[14674] <= 3'b000;
      memory_array[14675] <= 3'b000;
      memory_array[14676] <= 3'b000;
      memory_array[14677] <= 3'b101;
      memory_array[14678] <= 3'b101;
      memory_array[14679] <= 3'b111;
      memory_array[14680] <= 3'b111;
      memory_array[14681] <= 3'b111;
      memory_array[14682] <= 3'b101;
      memory_array[14683] <= 3'b101;
      memory_array[14684] <= 3'b101;
      memory_array[14685] <= 3'b101;
      memory_array[14686] <= 3'b101;
      memory_array[14687] <= 3'b101;
      memory_array[14688] <= 3'b000;
      memory_array[14689] <= 3'b000;
      memory_array[14690] <= 3'b000;
      memory_array[14691] <= 3'b000;
      memory_array[14692] <= 3'b000;
      memory_array[14693] <= 3'b000;
      memory_array[14694] <= 3'b000;
      memory_array[14695] <= 3'b000;
      memory_array[14696] <= 3'b000;
      memory_array[14697] <= 3'b101;
      memory_array[14698] <= 3'b101;
      memory_array[14699] <= 3'b101;
      memory_array[14700] <= 3'b101;
      memory_array[14701] <= 3'b101;
      memory_array[14702] <= 3'b101;
      memory_array[14703] <= 3'b101;
      memory_array[14704] <= 3'b101;
      memory_array[14705] <= 3'b101;
      memory_array[14706] <= 3'b101;
      memory_array[14707] <= 3'b101;
      memory_array[14708] <= 3'b000;
      memory_array[14709] <= 3'b000;
      memory_array[14710] <= 3'b000;
      memory_array[14711] <= 3'b101;
      memory_array[14712] <= 3'b101;
      memory_array[14713] <= 3'b000;
      memory_array[14714] <= 3'b000;
      memory_array[14715] <= 3'b101;
      memory_array[14716] <= 3'b101;
      memory_array[14717] <= 3'b000;
      memory_array[14718] <= 3'b000;
      memory_array[14719] <= 3'b000;
      memory_array[14720] <= 3'b101;
      memory_array[14721] <= 3'b101;
      memory_array[14722] <= 3'b101;
      memory_array[14723] <= 3'b101;
      memory_array[14724] <= 3'b000;
      memory_array[14725] <= 3'b000;
      memory_array[14726] <= 3'b101;
      memory_array[14727] <= 3'b101;
      memory_array[14728] <= 3'b101;
      memory_array[14729] <= 3'b000;
      memory_array[14730] <= 3'b101;
      memory_array[14731] <= 3'b101;
      memory_array[14732] <= 3'b000;
      memory_array[14733] <= 3'b000;
      memory_array[14734] <= 3'b000;
      memory_array[14735] <= 3'b000;
      memory_array[14736] <= 3'b000;
      memory_array[14737] <= 3'b000;
      memory_array[14738] <= 3'b000;
      memory_array[14739] <= 3'b000;
      memory_array[14740] <= 3'b000;
      memory_array[14741] <= 3'b000;
      memory_array[14742] <= 3'b000;
      memory_array[14743] <= 3'b000;
      memory_array[14744] <= 3'b000;
      memory_array[14745] <= 3'b110;
      memory_array[14746] <= 3'b000;
      memory_array[14747] <= 3'b000;
      memory_array[14748] <= 3'b000;
      memory_array[14749] <= 3'b000;
      memory_array[14750] <= 3'b111;
      memory_array[14751] <= 3'b111;
      memory_array[14752] <= 3'b111;
      memory_array[14753] <= 3'b111;
      memory_array[14754] <= 3'b111;
      memory_array[14755] <= 3'b101;
      memory_array[14756] <= 3'b101;
      memory_array[14757] <= 3'b101;
      memory_array[14758] <= 3'b101;
      memory_array[14759] <= 3'b101;
      memory_array[14760] <= 3'b101;
      memory_array[14761] <= 3'b111;
      memory_array[14762] <= 3'b111;
      memory_array[14763] <= 3'b111;
      memory_array[14764] <= 3'b111;
      memory_array[14765] <= 3'b111;
      memory_array[14766] <= 3'b101;
      memory_array[14767] <= 3'b101;
      memory_array[14768] <= 3'b101;
      memory_array[14769] <= 3'b101;
      memory_array[14770] <= 3'b101;
      memory_array[14771] <= 3'b111;
      memory_array[14772] <= 3'b111;
      memory_array[14773] <= 3'b111;
      memory_array[14774] <= 3'b111;
      memory_array[14775] <= 3'b111;
      memory_array[14776] <= 3'b101;
      memory_array[14777] <= 3'b101;
      memory_array[14778] <= 3'b101;
      memory_array[14779] <= 3'b101;
      memory_array[14780] <= 3'b101;
      memory_array[14781] <= 3'b111;
      memory_array[14782] <= 3'b111;
      memory_array[14783] <= 3'b111;
      memory_array[14784] <= 3'b111;
      memory_array[14785] <= 3'b111;
      memory_array[14786] <= 3'b101;
      memory_array[14787] <= 3'b101;
      memory_array[14788] <= 3'b101;
      memory_array[14789] <= 3'b000;
      memory_array[14790] <= 3'b000;
      memory_array[14791] <= 3'b101;
      memory_array[14792] <= 3'b110;
      memory_array[14793] <= 3'b000;
      memory_array[14794] <= 3'b000;
      memory_array[14795] <= 3'b110;
      memory_array[14796] <= 3'b110;
      memory_array[14797] <= 3'b110;
      memory_array[14798] <= 3'b000;
      memory_array[14799] <= 3'b101;
      memory_array[14800] <= 3'b101;
      memory_array[14801] <= 3'b101;
      memory_array[14802] <= 3'b110;
      memory_array[14803] <= 3'b101;
      memory_array[14804] <= 3'b101;
      memory_array[14805] <= 3'b110;
      memory_array[14806] <= 3'b101;
      memory_array[14807] <= 3'b101;
      memory_array[14808] <= 3'b101;
      memory_array[14809] <= 3'b000;
      memory_array[14810] <= 3'b000;
      memory_array[14811] <= 3'b101;
      memory_array[14812] <= 3'b101;
      memory_array[14813] <= 3'b101;
      memory_array[14814] <= 3'b111;
      memory_array[14815] <= 3'b111;
      memory_array[14816] <= 3'b111;
      memory_array[14817] <= 3'b111;
      memory_array[14818] <= 3'b111;
      memory_array[14819] <= 3'b101;
      memory_array[14820] <= 3'b101;
      memory_array[14821] <= 3'b101;
      memory_array[14822] <= 3'b101;
      memory_array[14823] <= 3'b101;
      memory_array[14824] <= 3'b111;
      memory_array[14825] <= 3'b111;
      memory_array[14826] <= 3'b111;
      memory_array[14827] <= 3'b111;
      memory_array[14828] <= 3'b111;
      memory_array[14829] <= 3'b101;
      memory_array[14830] <= 3'b101;
      memory_array[14831] <= 3'b101;
      memory_array[14832] <= 3'b101;
      memory_array[14833] <= 3'b101;
      memory_array[14834] <= 3'b111;
      memory_array[14835] <= 3'b111;
      memory_array[14836] <= 3'b111;
      memory_array[14837] <= 3'b111;
      memory_array[14838] <= 3'b111;
      memory_array[14839] <= 3'b101;
      memory_array[14840] <= 3'b101;
      memory_array[14841] <= 3'b101;
      memory_array[14842] <= 3'b101;
      memory_array[14843] <= 3'b101;
      memory_array[14844] <= 3'b111;
      memory_array[14845] <= 3'b111;
      memory_array[14846] <= 3'b111;
      memory_array[14847] <= 3'b111;
      memory_array[14848] <= 3'b111;
      memory_array[14849] <= 3'b101;
      memory_array[14850] <= 3'b000;
      memory_array[14851] <= 3'b000;
      memory_array[14852] <= 3'b000;
      memory_array[14853] <= 3'b000;
      memory_array[14854] <= 3'b000;
      memory_array[14855] <= 3'b000;
      memory_array[14856] <= 3'b101;
      memory_array[14857] <= 3'b101;
      memory_array[14858] <= 3'b000;
      memory_array[14859] <= 3'b000;
      memory_array[14860] <= 3'b000;
      memory_array[14861] <= 3'b000;
      memory_array[14862] <= 3'b000;
      memory_array[14863] <= 3'b000;
      memory_array[14864] <= 3'b000;
      memory_array[14865] <= 3'b000;
      memory_array[14866] <= 3'b000;
      memory_array[14867] <= 3'b000;
      memory_array[14868] <= 3'b000;
      memory_array[14869] <= 3'b000;
      memory_array[14870] <= 3'b110;
      memory_array[14871] <= 3'b000;
      memory_array[14872] <= 3'b000;
      memory_array[14873] <= 3'b000;
      memory_array[14874] <= 3'b000;
      memory_array[14875] <= 3'b000;
      memory_array[14876] <= 3'b000;
      memory_array[14877] <= 3'b101;
      memory_array[14878] <= 3'b101;
      memory_array[14879] <= 3'b101;
      memory_array[14880] <= 3'b101;
      memory_array[14881] <= 3'b111;
      memory_array[14882] <= 3'b111;
      memory_array[14883] <= 3'b111;
      memory_array[14884] <= 3'b101;
      memory_array[14885] <= 3'b101;
      memory_array[14886] <= 3'b101;
      memory_array[14887] <= 3'b101;
      memory_array[14888] <= 3'b000;
      memory_array[14889] <= 3'b000;
      memory_array[14890] <= 3'b000;
      memory_array[14891] <= 3'b101;
      memory_array[14892] <= 3'b111;
      memory_array[14893] <= 3'b111;
      memory_array[14894] <= 3'b111;
      memory_array[14895] <= 3'b111;
      memory_array[14896] <= 3'b111;
      memory_array[14897] <= 3'b111;
      memory_array[14898] <= 3'b111;
      memory_array[14899] <= 3'b111;
      memory_array[14900] <= 3'b111;
      memory_array[14901] <= 3'b101;
      memory_array[14902] <= 3'b101;
      memory_array[14903] <= 3'b101;
      memory_array[14904] <= 3'b000;
      memory_array[14905] <= 3'b000;
      memory_array[14906] <= 3'b000;
      memory_array[14907] <= 3'b000;
      memory_array[14908] <= 3'b000;
      memory_array[14909] <= 3'b101;
      memory_array[14910] <= 3'b101;
      memory_array[14911] <= 3'b101;
      memory_array[14912] <= 3'b101;
      memory_array[14913] <= 3'b000;
      memory_array[14914] <= 3'b000;
      memory_array[14915] <= 3'b101;
      memory_array[14916] <= 3'b101;
      memory_array[14917] <= 3'b000;
      memory_array[14918] <= 3'b000;
      memory_array[14919] <= 3'b000;
      memory_array[14920] <= 3'b000;
      memory_array[14921] <= 3'b000;
      memory_array[14922] <= 3'b000;
      memory_array[14923] <= 3'b000;
      memory_array[14924] <= 3'b000;
      memory_array[14925] <= 3'b000;
      memory_array[14926] <= 3'b000;
      memory_array[14927] <= 3'b000;
      memory_array[14928] <= 3'b000;
      memory_array[14929] <= 3'b101;
      memory_array[14930] <= 3'b101;
      memory_array[14931] <= 3'b000;
      memory_array[14932] <= 3'b110;
      memory_array[14933] <= 3'b000;
      memory_array[14934] <= 3'b000;
      memory_array[14935] <= 3'b000;
      memory_array[14936] <= 3'b000;
      memory_array[14937] <= 3'b000;
      memory_array[14938] <= 3'b000;
      memory_array[14939] <= 3'b000;
      memory_array[14940] <= 3'b000;
      memory_array[14941] <= 3'b000;
      memory_array[14942] <= 3'b000;
      memory_array[14943] <= 3'b000;
      memory_array[14944] <= 3'b000;
      memory_array[14945] <= 3'b101;
      memory_array[14946] <= 3'b000;
      memory_array[14947] <= 3'b000;
      memory_array[14948] <= 3'b000;
      memory_array[14949] <= 3'b000;
      memory_array[14950] <= 3'b111;
      memory_array[14951] <= 3'b111;
      memory_array[14952] <= 3'b111;
      memory_array[14953] <= 3'b111;
      memory_array[14954] <= 3'b111;
      memory_array[14955] <= 3'b101;
      memory_array[14956] <= 3'b101;
      memory_array[14957] <= 3'b101;
      memory_array[14958] <= 3'b101;
      memory_array[14959] <= 3'b101;
      memory_array[14960] <= 3'b101;
      memory_array[14961] <= 3'b111;
      memory_array[14962] <= 3'b111;
      memory_array[14963] <= 3'b111;
      memory_array[14964] <= 3'b111;
      memory_array[14965] <= 3'b111;
      memory_array[14966] <= 3'b101;
      memory_array[14967] <= 3'b101;
      memory_array[14968] <= 3'b101;
      memory_array[14969] <= 3'b101;
      memory_array[14970] <= 3'b101;
      memory_array[14971] <= 3'b111;
      memory_array[14972] <= 3'b111;
      memory_array[14973] <= 3'b111;
      memory_array[14974] <= 3'b111;
      memory_array[14975] <= 3'b111;
      memory_array[14976] <= 3'b101;
      memory_array[14977] <= 3'b101;
      memory_array[14978] <= 3'b101;
      memory_array[14979] <= 3'b101;
      memory_array[14980] <= 3'b101;
      memory_array[14981] <= 3'b111;
      memory_array[14982] <= 3'b111;
      memory_array[14983] <= 3'b111;
      memory_array[14984] <= 3'b111;
      memory_array[14985] <= 3'b111;
      memory_array[14986] <= 3'b101;
      memory_array[14987] <= 3'b101;
      memory_array[14988] <= 3'b101;
      memory_array[14989] <= 3'b000;
      memory_array[14990] <= 3'b000;
      memory_array[14991] <= 3'b101;
      memory_array[14992] <= 3'b101;
      memory_array[14993] <= 3'b101;
      memory_array[14994] <= 3'b000;
      memory_array[14995] <= 3'b101;
      memory_array[14996] <= 3'b101;
      memory_array[14997] <= 3'b110;
      memory_array[14998] <= 3'b101;
      memory_array[14999] <= 3'b101;
      // memory_array[15000] <= 3'b101;
      // memory_array[15001] <= 3'b101;
      // memory_array[15002] <= 3'b101;
      // memory_array[15003] <= 3'b111;
      // memory_array[15004] <= 3'b111;
      // memory_array[15005] <= 3'b101;
      // memory_array[15006] <= 3'b101;
      // memory_array[15007] <= 3'b101;
      // memory_array[15008] <= 3'b101;
      // memory_array[15009] <= 3'b000;
      // memory_array[15010] <= 3'b000;
      // memory_array[15011] <= 3'b101;
      // memory_array[15012] <= 3'b101;
      // memory_array[15013] <= 3'b101;
      // memory_array[15014] <= 3'b111;
      // memory_array[15015] <= 3'b111;
      // memory_array[15016] <= 3'b111;
      // memory_array[15017] <= 3'b111;
      // memory_array[15018] <= 3'b111;
      // memory_array[15019] <= 3'b101;
      // memory_array[15020] <= 3'b101;
      // memory_array[15021] <= 3'b101;
      // memory_array[15022] <= 3'b101;
      // memory_array[15023] <= 3'b101;
      // memory_array[15024] <= 3'b111;
      // memory_array[15025] <= 3'b111;
      // memory_array[15026] <= 3'b111;
      // memory_array[15027] <= 3'b111;
      // memory_array[15028] <= 3'b111;
      // memory_array[15029] <= 3'b101;
      // memory_array[15030] <= 3'b101;
      // memory_array[15031] <= 3'b101;
      // memory_array[15032] <= 3'b101;
      // memory_array[15033] <= 3'b101;
      // memory_array[15034] <= 3'b111;
      // memory_array[15035] <= 3'b111;
      // memory_array[15036] <= 3'b111;
      // memory_array[15037] <= 3'b111;
      // memory_array[15038] <= 3'b111;
      // memory_array[15039] <= 3'b101;
      // memory_array[15040] <= 3'b101;
      // memory_array[15041] <= 3'b101;
      // memory_array[15042] <= 3'b101;
      // memory_array[15043] <= 3'b101;
      // memory_array[15044] <= 3'b111;
      // memory_array[15045] <= 3'b111;
      // memory_array[15046] <= 3'b111;
      // memory_array[15047] <= 3'b111;
      // memory_array[15048] <= 3'b111;
      // memory_array[15049] <= 3'b101;
      // memory_array[15050] <= 3'b000;
      // memory_array[15051] <= 3'b000;
      // memory_array[15052] <= 3'b000;
      // memory_array[15053] <= 3'b000;
      // memory_array[15054] <= 3'b000;
      // memory_array[15055] <= 3'b000;
      // memory_array[15056] <= 3'b000;
      // memory_array[15057] <= 3'b000;
      // memory_array[15058] <= 3'b000;
      // memory_array[15059] <= 3'b000;
      // memory_array[15060] <= 3'b000;
      // memory_array[15061] <= 3'b000;
      // memory_array[15062] <= 3'b000;
      // memory_array[15063] <= 3'b000;
      // memory_array[15064] <= 3'b000;
      // memory_array[15065] <= 3'b000;
      // memory_array[15066] <= 3'b000;
      // memory_array[15067] <= 3'b000;
      // memory_array[15068] <= 3'b110;
      // memory_array[15069] <= 3'b000;
      // memory_array[15070] <= 3'b000;
      // memory_array[15071] <= 3'b000;
      // memory_array[15072] <= 3'b000;
      // memory_array[15073] <= 3'b000;
      // memory_array[15074] <= 3'b000;
      // memory_array[15075] <= 3'b000;
      // memory_array[15076] <= 3'b000;
      // memory_array[15077] <= 3'b101;
      // memory_array[15078] <= 3'b101;
      // memory_array[15079] <= 3'b111;
      // memory_array[15080] <= 3'b101;
      // memory_array[15081] <= 3'b111;
      // memory_array[15082] <= 3'b101;
      // memory_array[15083] <= 3'b111;
      // memory_array[15084] <= 3'b111;
      // memory_array[15085] <= 3'b101;
      // memory_array[15086] <= 3'b101;
      // memory_array[15087] <= 3'b101;
      // memory_array[15088] <= 3'b101;
      // memory_array[15089] <= 3'b101;
      // memory_array[15090] <= 3'b111;
      // memory_array[15091] <= 3'b111;
      // memory_array[15092] <= 3'b111;
      // memory_array[15093] <= 3'b101;
      // memory_array[15094] <= 3'b101;
      // memory_array[15095] <= 3'b101;
      // memory_array[15096] <= 3'b111;
      // memory_array[15097] <= 3'b101;
      // memory_array[15098] <= 3'b101;
      // memory_array[15099] <= 3'b101;
      // memory_array[15100] <= 3'b101;
      // memory_array[15101] <= 3'b101;
      // memory_array[15102] <= 3'b101;
      // memory_array[15103] <= 3'b101;
      // memory_array[15104] <= 3'b101;
      // memory_array[15105] <= 3'b101;
      // memory_array[15106] <= 3'b000;
      // memory_array[15107] <= 3'b000;
      // memory_array[15108] <= 3'b101;
      // memory_array[15109] <= 3'b101;
      // memory_array[15110] <= 3'b000;
      // memory_array[15111] <= 3'b101;
      // memory_array[15112] <= 3'b101;
      // memory_array[15113] <= 3'b101;
      // memory_array[15114] <= 3'b101;
      // memory_array[15115] <= 3'b000;
      // memory_array[15116] <= 3'b000;
      // memory_array[15117] <= 3'b000;
      // memory_array[15118] <= 3'b000;
      // memory_array[15119] <= 3'b000;
      // memory_array[15120] <= 3'b000;
      // memory_array[15121] <= 3'b000;
      // memory_array[15122] <= 3'b000;
      // memory_array[15123] <= 3'b000;
      // memory_array[15124] <= 3'b000;
      // memory_array[15125] <= 3'b000;
      // memory_array[15126] <= 3'b000;
      // memory_array[15127] <= 3'b000;
      // memory_array[15128] <= 3'b000;
      // memory_array[15129] <= 3'b000;
      // memory_array[15130] <= 3'b000;
      // memory_array[15131] <= 3'b000;
      // memory_array[15132] <= 3'b000;
      // memory_array[15133] <= 3'b000;
      // memory_array[15134] <= 3'b000;
      // memory_array[15135] <= 3'b000;
      // memory_array[15136] <= 3'b000;
      // memory_array[15137] <= 3'b000;
      // memory_array[15138] <= 3'b000;
      // memory_array[15139] <= 3'b000;
      // memory_array[15140] <= 3'b000;
      // memory_array[15141] <= 3'b000;
      // memory_array[15142] <= 3'b000;
      // memory_array[15143] <= 3'b110;
      // memory_array[15144] <= 3'b101;
      // memory_array[15145] <= 3'b000;
      // memory_array[15146] <= 3'b000;
      // memory_array[15147] <= 3'b000;
      // memory_array[15148] <= 3'b000;
      // memory_array[15149] <= 3'b000;
      // memory_array[15150] <= 3'b111;
      // memory_array[15151] <= 3'b111;
      // memory_array[15152] <= 3'b111;
      // memory_array[15153] <= 3'b111;
      // memory_array[15154] <= 3'b111;
      // memory_array[15155] <= 3'b101;
      // memory_array[15156] <= 3'b101;
      // memory_array[15157] <= 3'b101;
      // memory_array[15158] <= 3'b101;
      // memory_array[15159] <= 3'b101;
      // memory_array[15160] <= 3'b101;
      // memory_array[15161] <= 3'b111;
      // memory_array[15162] <= 3'b111;
      // memory_array[15163] <= 3'b111;
      // memory_array[15164] <= 3'b111;
      // memory_array[15165] <= 3'b111;
      // memory_array[15166] <= 3'b101;
      // memory_array[15167] <= 3'b101;
      // memory_array[15168] <= 3'b101;
      // memory_array[15169] <= 3'b101;
      // memory_array[15170] <= 3'b101;
      // memory_array[15171] <= 3'b111;
      // memory_array[15172] <= 3'b111;
      // memory_array[15173] <= 3'b111;
      // memory_array[15174] <= 3'b111;
      // memory_array[15175] <= 3'b111;
      // memory_array[15176] <= 3'b101;
      // memory_array[15177] <= 3'b101;
      // memory_array[15178] <= 3'b101;
      // memory_array[15179] <= 3'b101;
      // memory_array[15180] <= 3'b101;
      // memory_array[15181] <= 3'b111;
      // memory_array[15182] <= 3'b111;
      // memory_array[15183] <= 3'b111;
      // memory_array[15184] <= 3'b111;
      // memory_array[15185] <= 3'b111;
      // memory_array[15186] <= 3'b101;
      // memory_array[15187] <= 3'b101;
      // memory_array[15188] <= 3'b101;
      // memory_array[15189] <= 3'b000;
      // memory_array[15190] <= 3'b000;
      // memory_array[15191] <= 3'b101;
      // memory_array[15192] <= 3'b101;
      // memory_array[15193] <= 3'b101;
      // memory_array[15194] <= 3'b101;
      // memory_array[15195] <= 3'b111;
      // memory_array[15196] <= 3'b111;
      // memory_array[15197] <= 3'b101;
      // memory_array[15198] <= 3'b101;
      // memory_array[15199] <= 3'b101;
      // memory_array[15200] <= 3'b101;
      // memory_array[15201] <= 3'b101;
      // memory_array[15202] <= 3'b101;
      // memory_array[15203] <= 3'b101;
      // memory_array[15204] <= 3'b101;
      // memory_array[15205] <= 3'b101;
      // memory_array[15206] <= 3'b101;
      // memory_array[15207] <= 3'b101;
      // memory_array[15208] <= 3'b101;
      // memory_array[15209] <= 3'b000;
      // memory_array[15210] <= 3'b000;
      // memory_array[15211] <= 3'b101;
      // memory_array[15212] <= 3'b101;
      // memory_array[15213] <= 3'b101;
      // memory_array[15214] <= 3'b111;
      // memory_array[15215] <= 3'b111;
      // memory_array[15216] <= 3'b111;
      // memory_array[15217] <= 3'b111;
      // memory_array[15218] <= 3'b111;
      // memory_array[15219] <= 3'b101;
      // memory_array[15220] <= 3'b101;
      // memory_array[15221] <= 3'b101;
      // memory_array[15222] <= 3'b101;
      // memory_array[15223] <= 3'b101;
      // memory_array[15224] <= 3'b111;
      // memory_array[15225] <= 3'b111;
      // memory_array[15226] <= 3'b111;
      // memory_array[15227] <= 3'b111;
      // memory_array[15228] <= 3'b111;
      // memory_array[15229] <= 3'b101;
      // memory_array[15230] <= 3'b101;
      // memory_array[15231] <= 3'b101;
      // memory_array[15232] <= 3'b101;
      // memory_array[15233] <= 3'b101;
      // memory_array[15234] <= 3'b111;
      // memory_array[15235] <= 3'b111;
      // memory_array[15236] <= 3'b111;
      // memory_array[15237] <= 3'b111;
      // memory_array[15238] <= 3'b111;
      // memory_array[15239] <= 3'b101;
      // memory_array[15240] <= 3'b101;
      // memory_array[15241] <= 3'b101;
      // memory_array[15242] <= 3'b101;
      // memory_array[15243] <= 3'b101;
      // memory_array[15244] <= 3'b111;
      // memory_array[15245] <= 3'b111;
      // memory_array[15246] <= 3'b111;
      // memory_array[15247] <= 3'b111;
      // memory_array[15248] <= 3'b111;
      // memory_array[15249] <= 3'b101;
      // memory_array[15250] <= 3'b000;
      // memory_array[15251] <= 3'b000;
      // memory_array[15252] <= 3'b000;
      // memory_array[15253] <= 3'b000;
      // memory_array[15254] <= 3'b000;
      // memory_array[15255] <= 3'b000;
      // memory_array[15256] <= 3'b101;
      // memory_array[15257] <= 3'b000;
      // memory_array[15258] <= 3'b000;
      // memory_array[15259] <= 3'b000;
      // memory_array[15260] <= 3'b101;
      // memory_array[15261] <= 3'b101;
      // memory_array[15262] <= 3'b101;
      // memory_array[15263] <= 3'b000;
      // memory_array[15264] <= 3'b000;
      // memory_array[15265] <= 3'b101;
      // memory_array[15266] <= 3'b000;
      // memory_array[15267] <= 3'b110;
      // memory_array[15268] <= 3'b000;
      // memory_array[15269] <= 3'b000;
      // memory_array[15270] <= 3'b000;
      // memory_array[15271] <= 3'b110;
      // memory_array[15272] <= 3'b110;
      // memory_array[15273] <= 3'b000;
      // memory_array[15274] <= 3'b000;
      // memory_array[15275] <= 3'b000;
      // memory_array[15276] <= 3'b000;
      // memory_array[15277] <= 3'b101;
      // memory_array[15278] <= 3'b000;
      // memory_array[15279] <= 3'b101;
      // memory_array[15280] <= 3'b101;
      // memory_array[15281] <= 3'b101;
      // memory_array[15282] <= 3'b111;
      // memory_array[15283] <= 3'b111;
      // memory_array[15284] <= 3'b101;
      // memory_array[15285] <= 3'b111;
      // memory_array[15286] <= 3'b101;
      // memory_array[15287] <= 3'b101;
      // memory_array[15288] <= 3'b111;
      // memory_array[15289] <= 3'b111;
      // memory_array[15290] <= 3'b111;
      // memory_array[15291] <= 3'b111;
      // memory_array[15292] <= 3'b111;
      // memory_array[15293] <= 3'b101;
      // memory_array[15294] <= 3'b101;
      // memory_array[15295] <= 3'b101;
      // memory_array[15296] <= 3'b101;
      // memory_array[15297] <= 3'b101;
      // memory_array[15298] <= 3'b101;
      // memory_array[15299] <= 3'b000;
      // memory_array[15300] <= 3'b101;
      // memory_array[15301] <= 3'b101;
      // memory_array[15302] <= 3'b101;
      // memory_array[15303] <= 3'b000;
      // memory_array[15304] <= 3'b000;
      // memory_array[15305] <= 3'b101;
      // memory_array[15306] <= 3'b101;
      // memory_array[15307] <= 3'b000;
      // memory_array[15308] <= 3'b000;
      // memory_array[15309] <= 3'b000;
      // memory_array[15310] <= 3'b101;
      // memory_array[15311] <= 3'b101;
      // memory_array[15312] <= 3'b101;
      // memory_array[15313] <= 3'b000;
      // memory_array[15314] <= 3'b000;
      // memory_array[15315] <= 3'b101;
      // memory_array[15316] <= 3'b000;
      // memory_array[15317] <= 3'b000;
      // memory_array[15318] <= 3'b000;
      // memory_array[15319] <= 3'b000;
      // memory_array[15320] <= 3'b101;
      // memory_array[15321] <= 3'b110;
      // memory_array[15322] <= 3'b110;
      // memory_array[15323] <= 3'b000;
      // memory_array[15324] <= 3'b000;
      // memory_array[15325] <= 3'b000;
      // memory_array[15326] <= 3'b000;
      // memory_array[15327] <= 3'b000;
      // memory_array[15328] <= 3'b000;
      // memory_array[15329] <= 3'b000;
      // memory_array[15330] <= 3'b000;
      // memory_array[15331] <= 3'b000;
      // memory_array[15332] <= 3'b000;
      // memory_array[15333] <= 3'b000;
      // memory_array[15334] <= 3'b000;
      // memory_array[15335] <= 3'b000;
      // memory_array[15336] <= 3'b000;
      // memory_array[15337] <= 3'b000;
      // memory_array[15338] <= 3'b000;
      // memory_array[15339] <= 3'b000;
      // memory_array[15340] <= 3'b000;
      // memory_array[15341] <= 3'b000;
      // memory_array[15342] <= 3'b110;
      // memory_array[15343] <= 3'b000;
      // memory_array[15344] <= 3'b000;
      // memory_array[15345] <= 3'b110;
      // memory_array[15346] <= 3'b000;
      // memory_array[15347] <= 3'b000;
      // memory_array[15348] <= 3'b000;
      // memory_array[15349] <= 3'b000;
      // memory_array[15350] <= 3'b111;
      // memory_array[15351] <= 3'b111;
      // memory_array[15352] <= 3'b111;
      // memory_array[15353] <= 3'b111;
      // memory_array[15354] <= 3'b111;
      // memory_array[15355] <= 3'b101;
      // memory_array[15356] <= 3'b101;
      // memory_array[15357] <= 3'b101;
      // memory_array[15358] <= 3'b101;
      // memory_array[15359] <= 3'b101;
      // memory_array[15360] <= 3'b101;
      // memory_array[15361] <= 3'b111;
      // memory_array[15362] <= 3'b111;
      // memory_array[15363] <= 3'b111;
      // memory_array[15364] <= 3'b111;
      // memory_array[15365] <= 3'b111;
      // memory_array[15366] <= 3'b101;
      // memory_array[15367] <= 3'b101;
      // memory_array[15368] <= 3'b101;
      // memory_array[15369] <= 3'b101;
      // memory_array[15370] <= 3'b101;
      // memory_array[15371] <= 3'b111;
      // memory_array[15372] <= 3'b111;
      // memory_array[15373] <= 3'b111;
      // memory_array[15374] <= 3'b111;
      // memory_array[15375] <= 3'b111;
      // memory_array[15376] <= 3'b101;
      // memory_array[15377] <= 3'b101;
      // memory_array[15378] <= 3'b101;
      // memory_array[15379] <= 3'b101;
      // memory_array[15380] <= 3'b101;
      // memory_array[15381] <= 3'b111;
      // memory_array[15382] <= 3'b111;
      // memory_array[15383] <= 3'b111;
      // memory_array[15384] <= 3'b111;
      // memory_array[15385] <= 3'b111;
      // memory_array[15386] <= 3'b101;
      // memory_array[15387] <= 3'b101;
      // memory_array[15388] <= 3'b101;
      // memory_array[15389] <= 3'b000;
      // memory_array[15390] <= 3'b000;
      // memory_array[15391] <= 3'b101;
      // memory_array[15392] <= 3'b101;
      // memory_array[15393] <= 3'b101;
      // memory_array[15394] <= 3'b101;
      // memory_array[15395] <= 3'b101;
      // memory_array[15396] <= 3'b101;
      // memory_array[15397] <= 3'b101;
      // memory_array[15398] <= 3'b101;
      // memory_array[15399] <= 3'b101;
      // memory_array[15400] <= 3'b101;
      // memory_array[15401] <= 3'b101;
      // memory_array[15402] <= 3'b101;
      // memory_array[15403] <= 3'b101;
      // memory_array[15404] <= 3'b101;
      // memory_array[15405] <= 3'b101;
      // memory_array[15406] <= 3'b101;
      // memory_array[15407] <= 3'b101;
      // memory_array[15408] <= 3'b101;
      // memory_array[15409] <= 3'b000;
      // memory_array[15410] <= 3'b000;
      // memory_array[15411] <= 3'b000;
      // memory_array[15412] <= 3'b000;
      // memory_array[15413] <= 3'b000;
      // memory_array[15414] <= 3'b000;
      // memory_array[15415] <= 3'b000;
      // memory_array[15416] <= 3'b000;
      // memory_array[15417] <= 3'b000;
      // memory_array[15418] <= 3'b000;
      // memory_array[15419] <= 3'b000;
      // memory_array[15420] <= 3'b000;
      // memory_array[15421] <= 3'b000;
      // memory_array[15422] <= 3'b000;
      // memory_array[15423] <= 3'b000;
      // memory_array[15424] <= 3'b000;
      // memory_array[15425] <= 3'b000;
      // memory_array[15426] <= 3'b000;
      // memory_array[15427] <= 3'b000;
      // memory_array[15428] <= 3'b000;
      // memory_array[15429] <= 3'b000;
      // memory_array[15430] <= 3'b000;
      // memory_array[15431] <= 3'b000;
      // memory_array[15432] <= 3'b000;
      // memory_array[15433] <= 3'b000;
      // memory_array[15434] <= 3'b000;
      // memory_array[15435] <= 3'b000;
      // memory_array[15436] <= 3'b000;
      // memory_array[15437] <= 3'b000;
      // memory_array[15438] <= 3'b000;
      // memory_array[15439] <= 3'b000;
      // memory_array[15440] <= 3'b000;
      // memory_array[15441] <= 3'b000;
      // memory_array[15442] <= 3'b000;
      // memory_array[15443] <= 3'b000;
      // memory_array[15444] <= 3'b111;
      // memory_array[15445] <= 3'b111;
      // memory_array[15446] <= 3'b111;
      // memory_array[15447] <= 3'b111;
      // memory_array[15448] <= 3'b111;
      // memory_array[15449] <= 3'b101;
      // memory_array[15450] <= 3'b000;
      // memory_array[15451] <= 3'b000;
      // memory_array[15452] <= 3'b000;
      // memory_array[15453] <= 3'b000;
      // memory_array[15454] <= 3'b000;
      // memory_array[15455] <= 3'b000;
      // memory_array[15456] <= 3'b000;
      // memory_array[15457] <= 3'b110;
      // memory_array[15458] <= 3'b000;
      // memory_array[15459] <= 3'b000;
      // memory_array[15460] <= 3'b000;
      // memory_array[15461] <= 3'b101;
      // memory_array[15462] <= 3'b000;
      // memory_array[15463] <= 3'b000;
      // memory_array[15464] <= 3'b000;
      // memory_array[15465] <= 3'b101;
      // memory_array[15466] <= 3'b000;
      // memory_array[15467] <= 3'b000;
      // memory_array[15468] <= 3'b000;
      // memory_array[15469] <= 3'b000;
      // memory_array[15470] <= 3'b000;
      // memory_array[15471] <= 3'b110;
      // memory_array[15472] <= 3'b110;
      // memory_array[15473] <= 3'b000;
      // memory_array[15474] <= 3'b000;
      // memory_array[15475] <= 3'b000;
      // memory_array[15476] <= 3'b000;
      // memory_array[15477] <= 3'b000;
      // memory_array[15478] <= 3'b000;
      // memory_array[15479] <= 3'b101;
      // memory_array[15480] <= 3'b101;
      // memory_array[15481] <= 3'b101;
      // memory_array[15482] <= 3'b101;
      // memory_array[15483] <= 3'b111;
      // memory_array[15484] <= 3'b101;
      // memory_array[15485] <= 3'b101;
      // memory_array[15486] <= 3'b101;
      // memory_array[15487] <= 3'b101;
      // memory_array[15488] <= 3'b101;
      // memory_array[15489] <= 3'b101;
      // memory_array[15490] <= 3'b101;
      // memory_array[15491] <= 3'b101;
      // memory_array[15492] <= 3'b101;
      // memory_array[15493] <= 3'b101;
      // memory_array[15494] <= 3'b101;
      // memory_array[15495] <= 3'b101;
      // memory_array[15496] <= 3'b101;
      // memory_array[15497] <= 3'b101;
      // memory_array[15498] <= 3'b101;
      // memory_array[15499] <= 3'b101;
      // memory_array[15500] <= 3'b101;
      // memory_array[15501] <= 3'b101;
      // memory_array[15502] <= 3'b101;
      // memory_array[15503] <= 3'b000;
      // memory_array[15504] <= 3'b000;
      // memory_array[15505] <= 3'b101;
      // memory_array[15506] <= 3'b101;
      // memory_array[15507] <= 3'b101;
      // memory_array[15508] <= 3'b000;
      // memory_array[15509] <= 3'b000;
      // memory_array[15510] <= 3'b101;
      // memory_array[15511] <= 3'b101;
      // memory_array[15512] <= 3'b101;
      // memory_array[15513] <= 3'b000;
      // memory_array[15514] <= 3'b000;
      // memory_array[15515] <= 3'b101;
      // memory_array[15516] <= 3'b000;
      // memory_array[15517] <= 3'b101;
      // memory_array[15518] <= 3'b000;
      // memory_array[15519] <= 3'b000;
      // memory_array[15520] <= 3'b101;
      // memory_array[15521] <= 3'b101;
      // memory_array[15522] <= 3'b000;
      // memory_array[15523] <= 3'b000;
      // memory_array[15524] <= 3'b000;
      // memory_array[15525] <= 3'b000;
      // memory_array[15526] <= 3'b000;
      // memory_array[15527] <= 3'b101;
      // memory_array[15528] <= 3'b000;
      // memory_array[15529] <= 3'b000;
      // memory_array[15530] <= 3'b000;
      // memory_array[15531] <= 3'b000;
      // memory_array[15532] <= 3'b000;
      // memory_array[15533] <= 3'b000;
      // memory_array[15534] <= 3'b000;
      // memory_array[15535] <= 3'b000;
      // memory_array[15536] <= 3'b000;
      // memory_array[15537] <= 3'b000;
      // memory_array[15538] <= 3'b000;
      // memory_array[15539] <= 3'b000;
      // memory_array[15540] <= 3'b000;
      // memory_array[15541] <= 3'b000;
      // memory_array[15542] <= 3'b000;
      // memory_array[15543] <= 3'b000;
      // memory_array[15544] <= 3'b000;
      // memory_array[15545] <= 3'b000;
      // memory_array[15546] <= 3'b000;
      // memory_array[15547] <= 3'b000;
      // memory_array[15548] <= 3'b000;
      // memory_array[15549] <= 3'b000;
      // memory_array[15550] <= 3'b111;
      // memory_array[15551] <= 3'b111;
      // memory_array[15552] <= 3'b111;
      // memory_array[15553] <= 3'b111;
      // memory_array[15554] <= 3'b111;
      // memory_array[15555] <= 3'b101;
      // memory_array[15556] <= 3'b000;
      // memory_array[15557] <= 3'b000;
      // memory_array[15558] <= 3'b000;
      // memory_array[15559] <= 3'b000;
      // memory_array[15560] <= 3'b000;
      // memory_array[15561] <= 3'b000;
      // memory_array[15562] <= 3'b000;
      // memory_array[15563] <= 3'b000;
      // memory_array[15564] <= 3'b000;
      // memory_array[15565] <= 3'b000;
      // memory_array[15566] <= 3'b000;
      // memory_array[15567] <= 3'b000;
      // memory_array[15568] <= 3'b000;
      // memory_array[15569] <= 3'b000;
      // memory_array[15570] <= 3'b000;
      // memory_array[15571] <= 3'b000;
      // memory_array[15572] <= 3'b000;
      // memory_array[15573] <= 3'b000;
      // memory_array[15574] <= 3'b000;
      // memory_array[15575] <= 3'b000;
      // memory_array[15576] <= 3'b000;
      // memory_array[15577] <= 3'b000;
      // memory_array[15578] <= 3'b000;
      // memory_array[15579] <= 3'b000;
      // memory_array[15580] <= 3'b000;
      // memory_array[15581] <= 3'b000;
      // memory_array[15582] <= 3'b000;
      // memory_array[15583] <= 3'b000;
      // memory_array[15584] <= 3'b000;
      // memory_array[15585] <= 3'b000;
      // memory_array[15586] <= 3'b000;
      // memory_array[15587] <= 3'b000;
      // memory_array[15588] <= 3'b000;
      // memory_array[15589] <= 3'b000;
      // memory_array[15590] <= 3'b000;
      // memory_array[15591] <= 3'b101;
      // memory_array[15592] <= 3'b101;
      // memory_array[15593] <= 3'b101;
      // memory_array[15594] <= 3'b101;
      // memory_array[15595] <= 3'b101;
      // memory_array[15596] <= 3'b101;
      // memory_array[15597] <= 3'b101;
      // memory_array[15598] <= 3'b101;
      // memory_array[15599] <= 3'b101;
      // memory_array[15600] <= 3'b101;
      // memory_array[15601] <= 3'b101;
      // memory_array[15602] <= 3'b101;
      // memory_array[15603] <= 3'b111;
      // memory_array[15604] <= 3'b111;
      // memory_array[15605] <= 3'b101;
      // memory_array[15606] <= 3'b101;
      // memory_array[15607] <= 3'b101;
      // memory_array[15608] <= 3'b101;
      // memory_array[15609] <= 3'b000;
      // memory_array[15610] <= 3'b000;
      // memory_array[15611] <= 3'b110;
      // memory_array[15612] <= 3'b000;
      // memory_array[15613] <= 3'b110;
      // memory_array[15614] <= 3'b110;
      // memory_array[15615] <= 3'b000;
      // memory_array[15616] <= 3'b111;
      // memory_array[15617] <= 3'b000;
      // memory_array[15618] <= 3'b110;
      // memory_array[15619] <= 3'b110;
      // memory_array[15620] <= 3'b000;
      // memory_array[15621] <= 3'b111;
      // memory_array[15622] <= 3'b000;
      // memory_array[15623] <= 3'b110;
      // memory_array[15624] <= 3'b110;
      // memory_array[15625] <= 3'b000;
      // memory_array[15626] <= 3'b111;
      // memory_array[15627] <= 3'b000;
      // memory_array[15628] <= 3'b110;
      // memory_array[15629] <= 3'b110;
      // memory_array[15630] <= 3'b000;
      // memory_array[15631] <= 3'b111;
      // memory_array[15632] <= 3'b000;
      // memory_array[15633] <= 3'b110;
      // memory_array[15634] <= 3'b110;
      // memory_array[15635] <= 3'b000;
      // memory_array[15636] <= 3'b111;
      // memory_array[15637] <= 3'b000;
      // memory_array[15638] <= 3'b110;
      // memory_array[15639] <= 3'b110;
      // memory_array[15640] <= 3'b000;
      // memory_array[15641] <= 3'b110;
      // memory_array[15642] <= 3'b000;
      // memory_array[15643] <= 3'b110;
      // memory_array[15644] <= 3'b111;
      // memory_array[15645] <= 3'b111;
      // memory_array[15646] <= 3'b111;
      // memory_array[15647] <= 3'b111;
      // memory_array[15648] <= 3'b111;
      // memory_array[15649] <= 3'b101;
      // memory_array[15650] <= 3'b000;
      // memory_array[15651] <= 3'b000;
      // memory_array[15652] <= 3'b000;
      // memory_array[15653] <= 3'b000;
      // memory_array[15654] <= 3'b000;
      // memory_array[15655] <= 3'b000;
      // memory_array[15656] <= 3'b000;
      // memory_array[15657] <= 3'b000;
      // memory_array[15658] <= 3'b110;
      // memory_array[15659] <= 3'b000;
      // memory_array[15660] <= 3'b000;
      // memory_array[15661] <= 3'b000;
      // memory_array[15662] <= 3'b000;
      // memory_array[15663] <= 3'b101;
      // memory_array[15664] <= 3'b000;
      // memory_array[15665] <= 3'b000;
      // memory_array[15666] <= 3'b000;
      // memory_array[15667] <= 3'b000;
      // memory_array[15668] <= 3'b000;
      // memory_array[15669] <= 3'b000;
      // memory_array[15670] <= 3'b000;
      // memory_array[15671] <= 3'b000;
      // memory_array[15672] <= 3'b000;
      // memory_array[15673] <= 3'b000;
      // memory_array[15674] <= 3'b000;
      // memory_array[15675] <= 3'b000;
      // memory_array[15676] <= 3'b000;
      // memory_array[15677] <= 3'b000;
      // memory_array[15678] <= 3'b000;
      // memory_array[15679] <= 3'b101;
      // memory_array[15680] <= 3'b000;
      // memory_array[15681] <= 3'b101;
      // memory_array[15682] <= 3'b101;
      // memory_array[15683] <= 3'b101;
      // memory_array[15684] <= 3'b101;
      // memory_array[15685] <= 3'b101;
      // memory_array[15686] <= 3'b101;
      // memory_array[15687] <= 3'b101;
      // memory_array[15688] <= 3'b101;
      // memory_array[15689] <= 3'b101;
      // memory_array[15690] <= 3'b101;
      // memory_array[15691] <= 3'b101;
      // memory_array[15692] <= 3'b101;
      // memory_array[15693] <= 3'b101;
      // memory_array[15694] <= 3'b101;
      // memory_array[15695] <= 3'b101;
      // memory_array[15696] <= 3'b101;
      // memory_array[15697] <= 3'b000;
      // memory_array[15698] <= 3'b101;
      // memory_array[15699] <= 3'b101;
      // memory_array[15700] <= 3'b000;
      // memory_array[15701] <= 3'b000;
      // memory_array[15702] <= 3'b000;
      // memory_array[15703] <= 3'b101;
      // memory_array[15704] <= 3'b101;
      // memory_array[15705] <= 3'b000;
      // memory_array[15706] <= 3'b000;
      // memory_array[15707] <= 3'b000;
      // memory_array[15708] <= 3'b101;
      // memory_array[15709] <= 3'b101;
      // memory_array[15710] <= 3'b000;
      // memory_array[15711] <= 3'b000;
      // memory_array[15712] <= 3'b000;
      // memory_array[15713] <= 3'b101;
      // memory_array[15714] <= 3'b101;
      // memory_array[15715] <= 3'b000;
      // memory_array[15716] <= 3'b000;
      // memory_array[15717] <= 3'b000;
      // memory_array[15718] <= 3'b000;
      // memory_array[15719] <= 3'b000;
      // memory_array[15720] <= 3'b000;
      // memory_array[15721] <= 3'b000;
      // memory_array[15722] <= 3'b000;
      // memory_array[15723] <= 3'b000;
      // memory_array[15724] <= 3'b000;
      // memory_array[15725] <= 3'b000;
      // memory_array[15726] <= 3'b000;
      // memory_array[15727] <= 3'b000;
      // memory_array[15728] <= 3'b000;
      // memory_array[15729] <= 3'b000;
      // memory_array[15730] <= 3'b000;
      // memory_array[15731] <= 3'b000;
      // memory_array[15732] <= 3'b000;
      // memory_array[15733] <= 3'b000;
      // memory_array[15734] <= 3'b000;
      // memory_array[15735] <= 3'b000;
      // memory_array[15736] <= 3'b000;
      // memory_array[15737] <= 3'b000;
      // memory_array[15738] <= 3'b000;
      // memory_array[15739] <= 3'b000;
      // memory_array[15740] <= 3'b000;
      // memory_array[15741] <= 3'b000;
      // memory_array[15742] <= 3'b000;
      // memory_array[15743] <= 3'b000;
      // memory_array[15744] <= 3'b000;
      // memory_array[15745] <= 3'b000;
      // memory_array[15746] <= 3'b000;
      // memory_array[15747] <= 3'b000;
      // memory_array[15748] <= 3'b000;
      // memory_array[15749] <= 3'b000;
      // memory_array[15750] <= 3'b111;
      // memory_array[15751] <= 3'b111;
      // memory_array[15752] <= 3'b111;
      // memory_array[15753] <= 3'b111;
      // memory_array[15754] <= 3'b111;
      // memory_array[15755] <= 3'b101;
      // memory_array[15756] <= 3'b000;
      // memory_array[15757] <= 3'b110;
      // memory_array[15758] <= 3'b110;
      // memory_array[15759] <= 3'b110;
      // memory_array[15760] <= 3'b110;
      // memory_array[15761] <= 3'b000;
      // memory_array[15762] <= 3'b111;
      // memory_array[15763] <= 3'b110;
      // memory_array[15764] <= 3'b110;
      // memory_array[15765] <= 3'b110;
      // memory_array[15766] <= 3'b000;
      // memory_array[15767] <= 3'b111;
      // memory_array[15768] <= 3'b110;
      // memory_array[15769] <= 3'b110;
      // memory_array[15770] <= 3'b111;
      // memory_array[15771] <= 3'b000;
      // memory_array[15772] <= 3'b111;
      // memory_array[15773] <= 3'b110;
      // memory_array[15774] <= 3'b110;
      // memory_array[15775] <= 3'b111;
      // memory_array[15776] <= 3'b000;
      // memory_array[15777] <= 3'b111;
      // memory_array[15778] <= 3'b110;
      // memory_array[15779] <= 3'b110;
      // memory_array[15780] <= 3'b111;
      // memory_array[15781] <= 3'b000;
      // memory_array[15782] <= 3'b111;
      // memory_array[15783] <= 3'b110;
      // memory_array[15784] <= 3'b110;
      // memory_array[15785] <= 3'b111;
      // memory_array[15786] <= 3'b000;
      // memory_array[15787] <= 3'b110;
      // memory_array[15788] <= 3'b110;
      // memory_array[15789] <= 3'b000;
      // memory_array[15790] <= 3'b000;
      // memory_array[15791] <= 3'b101;
      // memory_array[15792] <= 3'b101;
      // memory_array[15793] <= 3'b101;
      // memory_array[15794] <= 3'b101;
      // memory_array[15795] <= 3'b111;
      // memory_array[15796] <= 3'b111;
      // memory_array[15797] <= 3'b101;
      // memory_array[15798] <= 3'b101;
      // memory_array[15799] <= 3'b101;
      // memory_array[15800] <= 3'b101;
      // memory_array[15801] <= 3'b000;
      // memory_array[15802] <= 3'b000;
      // memory_array[15803] <= 3'b110;
      // memory_array[15804] <= 3'b110;
      // memory_array[15805] <= 3'b000;
      // memory_array[15806] <= 3'b000;
      // memory_array[15807] <= 3'b101;
      // memory_array[15808] <= 3'b101;
      // memory_array[15809] <= 3'b000;
      // memory_array[15810] <= 3'b000;
      // memory_array[15811] <= 3'b000;
      // memory_array[15812] <= 3'b000;
      // memory_array[15813] <= 3'b000;
      // memory_array[15814] <= 3'b000;
      // memory_array[15815] <= 3'b000;
      // memory_array[15816] <= 3'b000;
      // memory_array[15817] <= 3'b000;
      // memory_array[15818] <= 3'b000;
      // memory_array[15819] <= 3'b000;
      // memory_array[15820] <= 3'b000;
      // memory_array[15821] <= 3'b000;
      // memory_array[15822] <= 3'b000;
      // memory_array[15823] <= 3'b000;
      // memory_array[15824] <= 3'b000;
      // memory_array[15825] <= 3'b000;
      // memory_array[15826] <= 3'b000;
      // memory_array[15827] <= 3'b000;
      // memory_array[15828] <= 3'b000;
      // memory_array[15829] <= 3'b000;
      // memory_array[15830] <= 3'b000;
      // memory_array[15831] <= 3'b000;
      // memory_array[15832] <= 3'b000;
      // memory_array[15833] <= 3'b000;
      // memory_array[15834] <= 3'b000;
      // memory_array[15835] <= 3'b000;
      // memory_array[15836] <= 3'b000;
      // memory_array[15837] <= 3'b000;
      // memory_array[15838] <= 3'b000;
      // memory_array[15839] <= 3'b000;
      // memory_array[15840] <= 3'b000;
      // memory_array[15841] <= 3'b000;
      // memory_array[15842] <= 3'b000;
      // memory_array[15843] <= 3'b000;
      // memory_array[15844] <= 3'b110;
      // memory_array[15845] <= 3'b000;
      // memory_array[15846] <= 3'b000;
      // memory_array[15847] <= 3'b000;
      // memory_array[15848] <= 3'b000;
      // memory_array[15849] <= 3'b000;
      // memory_array[15850] <= 3'b000;
      // memory_array[15851] <= 3'b000;
      // memory_array[15852] <= 3'b000;
      // memory_array[15853] <= 3'b000;
      // memory_array[15854] <= 3'b000;
      // memory_array[15855] <= 3'b000;
      // memory_array[15856] <= 3'b000;
      // memory_array[15857] <= 3'b000;
      // memory_array[15858] <= 3'b000;
      // memory_array[15859] <= 3'b110;
      // memory_array[15860] <= 3'b000;
      // memory_array[15861] <= 3'b000;
      // memory_array[15862] <= 3'b000;
      // memory_array[15863] <= 3'b101;
      // memory_array[15864] <= 3'b000;
      // memory_array[15865] <= 3'b000;
      // memory_array[15866] <= 3'b000;
      // memory_array[15867] <= 3'b000;
      // memory_array[15868] <= 3'b000;
      // memory_array[15869] <= 3'b000;
      // memory_array[15870] <= 3'b000;
      // memory_array[15871] <= 3'b000;
      // memory_array[15872] <= 3'b000;
      // memory_array[15873] <= 3'b000;
      // memory_array[15874] <= 3'b000;
      // memory_array[15875] <= 3'b000;
      // memory_array[15876] <= 3'b000;
      // memory_array[15877] <= 3'b000;
      // memory_array[15878] <= 3'b000;
      // memory_array[15879] <= 3'b000;
      // memory_array[15880] <= 3'b000;
      // memory_array[15881] <= 3'b000;
      // memory_array[15882] <= 3'b000;
      // memory_array[15883] <= 3'b000;
      // memory_array[15884] <= 3'b000;
      // memory_array[15885] <= 3'b000;
      // memory_array[15886] <= 3'b000;
      // memory_array[15887] <= 3'b000;
      // memory_array[15888] <= 3'b000;
      // memory_array[15889] <= 3'b101;
      // memory_array[15890] <= 3'b000;
      // memory_array[15891] <= 3'b000;
      // memory_array[15892] <= 3'b000;
      // memory_array[15893] <= 3'b000;
      // memory_array[15894] <= 3'b000;
      // memory_array[15895] <= 3'b101;
      // memory_array[15896] <= 3'b101;
      // memory_array[15897] <= 3'b101;
      // memory_array[15898] <= 3'b101;
      // memory_array[15899] <= 3'b101;
      // memory_array[15900] <= 3'b000;
      // memory_array[15901] <= 3'b000;
      // memory_array[15902] <= 3'b000;
      // memory_array[15903] <= 3'b000;
      // memory_array[15904] <= 3'b000;
      // memory_array[15905] <= 3'b000;
      // memory_array[15906] <= 3'b000;
      // memory_array[15907] <= 3'b000;
      // memory_array[15908] <= 3'b101;
      // memory_array[15909] <= 3'b000;
      // memory_array[15910] <= 3'b000;
      // memory_array[15911] <= 3'b000;
      // memory_array[15912] <= 3'b000;
      // memory_array[15913] <= 3'b101;
      // memory_array[15914] <= 3'b000;
      // memory_array[15915] <= 3'b000;
      // memory_array[15916] <= 3'b000;
      // memory_array[15917] <= 3'b000;
      // memory_array[15918] <= 3'b000;
      // memory_array[15919] <= 3'b000;
      // memory_array[15920] <= 3'b000;
      // memory_array[15921] <= 3'b000;
      // memory_array[15922] <= 3'b000;
      // memory_array[15923] <= 3'b000;
      // memory_array[15924] <= 3'b000;
      // memory_array[15925] <= 3'b000;
      // memory_array[15926] <= 3'b000;
      // memory_array[15927] <= 3'b000;
      // memory_array[15928] <= 3'b000;
      // memory_array[15929] <= 3'b000;
      // memory_array[15930] <= 3'b000;
      // memory_array[15931] <= 3'b000;
      // memory_array[15932] <= 3'b000;
      // memory_array[15933] <= 3'b000;
      // memory_array[15934] <= 3'b101;
      // memory_array[15935] <= 3'b000;
      // memory_array[15936] <= 3'b000;
      // memory_array[15937] <= 3'b000;
      // memory_array[15938] <= 3'b000;
      // memory_array[15939] <= 3'b000;
      // memory_array[15940] <= 3'b000;
      // memory_array[15941] <= 3'b000;
      // memory_array[15942] <= 3'b000;
      // memory_array[15943] <= 3'b000;
      // memory_array[15944] <= 3'b000;
      // memory_array[15945] <= 3'b000;
      // memory_array[15946] <= 3'b000;
      // memory_array[15947] <= 3'b000;
      // memory_array[15948] <= 3'b000;
      // memory_array[15949] <= 3'b000;
      // memory_array[15950] <= 3'b110;
      // memory_array[15951] <= 3'b000;
      // memory_array[15952] <= 3'b000;
      // memory_array[15953] <= 3'b000;
      // memory_array[15954] <= 3'b000;
      // memory_array[15955] <= 3'b000;
      // memory_array[15956] <= 3'b000;
      // memory_array[15957] <= 3'b000;
      // memory_array[15958] <= 3'b000;
      // memory_array[15959] <= 3'b000;
      // memory_array[15960] <= 3'b000;
      // memory_array[15961] <= 3'b000;
      // memory_array[15962] <= 3'b000;
      // memory_array[15963] <= 3'b000;
      // memory_array[15964] <= 3'b000;
      // memory_array[15965] <= 3'b000;
      // memory_array[15966] <= 3'b000;
      // memory_array[15967] <= 3'b000;
      // memory_array[15968] <= 3'b000;
      // memory_array[15969] <= 3'b000;
      // memory_array[15970] <= 3'b000;
      // memory_array[15971] <= 3'b000;
      // memory_array[15972] <= 3'b000;
      // memory_array[15973] <= 3'b000;
      // memory_array[15974] <= 3'b000;
      // memory_array[15975] <= 3'b000;
      // memory_array[15976] <= 3'b000;
      // memory_array[15977] <= 3'b000;
      // memory_array[15978] <= 3'b000;
      // memory_array[15979] <= 3'b000;
      // memory_array[15980] <= 3'b000;
      // memory_array[15981] <= 3'b000;
      // memory_array[15982] <= 3'b000;
      // memory_array[15983] <= 3'b000;
      // memory_array[15984] <= 3'b000;
      // memory_array[15985] <= 3'b000;
      // memory_array[15986] <= 3'b000;
      // memory_array[15987] <= 3'b000;
      // memory_array[15988] <= 3'b000;
      // memory_array[15989] <= 3'b000;
      // memory_array[15990] <= 3'b000;
      // memory_array[15991] <= 3'b101;
      // memory_array[15992] <= 3'b101;
      // memory_array[15993] <= 3'b110;
      // memory_array[15994] <= 3'b110;
      // memory_array[15995] <= 3'b000;
      // memory_array[15996] <= 3'b000;
      // memory_array[15997] <= 3'b000;
      // memory_array[15998] <= 3'b110;
      // memory_array[15999] <= 3'b101;
      // memory_array[16000] <= 3'b101;
      // memory_array[16001] <= 3'b000;
      // memory_array[16002] <= 3'b000;
      // memory_array[16003] <= 3'b110;
      // memory_array[16004] <= 3'b110;
      // memory_array[16005] <= 3'b000;
      // memory_array[16006] <= 3'b000;
      // memory_array[16007] <= 3'b101;
      // memory_array[16008] <= 3'b101;
      // memory_array[16009] <= 3'b000;
      // memory_array[16010] <= 3'b000;
      // memory_array[16011] <= 3'b000;
      // memory_array[16012] <= 3'b000;
      // memory_array[16013] <= 3'b000;
      // memory_array[16014] <= 3'b000;
      // memory_array[16015] <= 3'b000;
      // memory_array[16016] <= 3'b000;
      // memory_array[16017] <= 3'b000;
      // memory_array[16018] <= 3'b000;
      // memory_array[16019] <= 3'b000;
      // memory_array[16020] <= 3'b000;
      // memory_array[16021] <= 3'b000;
      // memory_array[16022] <= 3'b000;
      // memory_array[16023] <= 3'b000;
      // memory_array[16024] <= 3'b000;
      // memory_array[16025] <= 3'b000;
      // memory_array[16026] <= 3'b000;
      // memory_array[16027] <= 3'b000;
      // memory_array[16028] <= 3'b000;
      // memory_array[16029] <= 3'b000;
      // memory_array[16030] <= 3'b000;
      // memory_array[16031] <= 3'b000;
      // memory_array[16032] <= 3'b000;
      // memory_array[16033] <= 3'b000;
      // memory_array[16034] <= 3'b000;
      // memory_array[16035] <= 3'b000;
      // memory_array[16036] <= 3'b000;
      // memory_array[16037] <= 3'b000;
      // memory_array[16038] <= 3'b000;
      // memory_array[16039] <= 3'b000;
      // memory_array[16040] <= 3'b000;
      // memory_array[16041] <= 3'b000;
      // memory_array[16042] <= 3'b000;
      // memory_array[16043] <= 3'b000;
      // memory_array[16044] <= 3'b110;
      // memory_array[16045] <= 3'b000;
      // memory_array[16046] <= 3'b000;
      // memory_array[16047] <= 3'b000;
      // memory_array[16048] <= 3'b000;
      // memory_array[16049] <= 3'b000;
      // memory_array[16050] <= 3'b000;
      // memory_array[16051] <= 3'b000;
      // memory_array[16052] <= 3'b000;
      // memory_array[16053] <= 3'b000;
      // memory_array[16054] <= 3'b000;
      // memory_array[16055] <= 3'b000;
      // memory_array[16056] <= 3'b000;
      // memory_array[16057] <= 3'b000;
      // memory_array[16058] <= 3'b000;
      // memory_array[16059] <= 3'b110;
      // memory_array[16060] <= 3'b000;
      // memory_array[16061] <= 3'b000;
      // memory_array[16062] <= 3'b000;
      // memory_array[16063] <= 3'b101;
      // memory_array[16064] <= 3'b000;
      // memory_array[16065] <= 3'b000;
      // memory_array[16066] <= 3'b000;
      // memory_array[16067] <= 3'b000;
      // memory_array[16068] <= 3'b000;
      // memory_array[16069] <= 3'b000;
      // memory_array[16070] <= 3'b000;
      // memory_array[16071] <= 3'b000;
      // memory_array[16072] <= 3'b000;
      // memory_array[16073] <= 3'b000;
      // memory_array[16074] <= 3'b000;
      // memory_array[16075] <= 3'b000;
      // memory_array[16076] <= 3'b000;
      // memory_array[16077] <= 3'b000;
      // memory_array[16078] <= 3'b000;
      // memory_array[16079] <= 3'b000;
      // memory_array[16080] <= 3'b000;
      // memory_array[16081] <= 3'b000;
      // memory_array[16082] <= 3'b000;
      // memory_array[16083] <= 3'b000;
      // memory_array[16084] <= 3'b000;
      // memory_array[16085] <= 3'b000;
      // memory_array[16086] <= 3'b000;
      // memory_array[16087] <= 3'b000;
      // memory_array[16088] <= 3'b000;
      // memory_array[16089] <= 3'b101;
      // memory_array[16090] <= 3'b000;
      // memory_array[16091] <= 3'b000;
      // memory_array[16092] <= 3'b000;
      // memory_array[16093] <= 3'b000;
      // memory_array[16094] <= 3'b000;
      // memory_array[16095] <= 3'b101;
      // memory_array[16096] <= 3'b101;
      // memory_array[16097] <= 3'b101;
      // memory_array[16098] <= 3'b101;
      // memory_array[16099] <= 3'b101;
      // memory_array[16100] <= 3'b000;
      // memory_array[16101] <= 3'b000;
      // memory_array[16102] <= 3'b000;
      // memory_array[16103] <= 3'b000;
      // memory_array[16104] <= 3'b000;
      // memory_array[16105] <= 3'b000;
      // memory_array[16106] <= 3'b000;
      // memory_array[16107] <= 3'b000;
      // memory_array[16108] <= 3'b101;
      // memory_array[16109] <= 3'b000;
      // memory_array[16110] <= 3'b000;
      // memory_array[16111] <= 3'b000;
      // memory_array[16112] <= 3'b000;
      // memory_array[16113] <= 3'b101;
      // memory_array[16114] <= 3'b000;
      // memory_array[16115] <= 3'b000;
      // memory_array[16116] <= 3'b000;
      // memory_array[16117] <= 3'b000;
      // memory_array[16118] <= 3'b000;
      // memory_array[16119] <= 3'b000;
      // memory_array[16120] <= 3'b000;
      // memory_array[16121] <= 3'b000;
      // memory_array[16122] <= 3'b000;
      // memory_array[16123] <= 3'b000;
      // memory_array[16124] <= 3'b000;
      // memory_array[16125] <= 3'b000;
      // memory_array[16126] <= 3'b000;
      // memory_array[16127] <= 3'b000;
      // memory_array[16128] <= 3'b000;
      // memory_array[16129] <= 3'b000;
      // memory_array[16130] <= 3'b000;
      // memory_array[16131] <= 3'b000;
      // memory_array[16132] <= 3'b000;
      // memory_array[16133] <= 3'b000;
      // memory_array[16134] <= 3'b101;
      // memory_array[16135] <= 3'b000;
      // memory_array[16136] <= 3'b000;
      // memory_array[16137] <= 3'b000;
      // memory_array[16138] <= 3'b000;
      // memory_array[16139] <= 3'b000;
      // memory_array[16140] <= 3'b000;
      // memory_array[16141] <= 3'b000;
      // memory_array[16142] <= 3'b000;
      // memory_array[16143] <= 3'b000;
      // memory_array[16144] <= 3'b000;
      // memory_array[16145] <= 3'b000;
      // memory_array[16146] <= 3'b000;
      // memory_array[16147] <= 3'b000;
      // memory_array[16148] <= 3'b000;
      // memory_array[16149] <= 3'b000;
      // memory_array[16150] <= 3'b110;
      // memory_array[16151] <= 3'b000;
      // memory_array[16152] <= 3'b000;
      // memory_array[16153] <= 3'b000;
      // memory_array[16154] <= 3'b000;
      // memory_array[16155] <= 3'b000;
      // memory_array[16156] <= 3'b000;
      // memory_array[16157] <= 3'b000;
      // memory_array[16158] <= 3'b000;
      // memory_array[16159] <= 3'b000;
      // memory_array[16160] <= 3'b000;
      // memory_array[16161] <= 3'b000;
      // memory_array[16162] <= 3'b000;
      // memory_array[16163] <= 3'b000;
      // memory_array[16164] <= 3'b000;
      // memory_array[16165] <= 3'b000;
      // memory_array[16166] <= 3'b000;
      // memory_array[16167] <= 3'b000;
      // memory_array[16168] <= 3'b000;
      // memory_array[16169] <= 3'b000;
      // memory_array[16170] <= 3'b000;
      // memory_array[16171] <= 3'b000;
      // memory_array[16172] <= 3'b000;
      // memory_array[16173] <= 3'b000;
      // memory_array[16174] <= 3'b000;
      // memory_array[16175] <= 3'b000;
      // memory_array[16176] <= 3'b000;
      // memory_array[16177] <= 3'b000;
      // memory_array[16178] <= 3'b000;
      // memory_array[16179] <= 3'b000;
      // memory_array[16180] <= 3'b000;
      // memory_array[16181] <= 3'b000;
      // memory_array[16182] <= 3'b000;
      // memory_array[16183] <= 3'b000;
      // memory_array[16184] <= 3'b000;
      // memory_array[16185] <= 3'b000;
      // memory_array[16186] <= 3'b000;
      // memory_array[16187] <= 3'b000;
      // memory_array[16188] <= 3'b000;
      // memory_array[16189] <= 3'b000;
      // memory_array[16190] <= 3'b000;
      // memory_array[16191] <= 3'b101;
      // memory_array[16192] <= 3'b101;
      // memory_array[16193] <= 3'b110;
      // memory_array[16194] <= 3'b110;
      // memory_array[16195] <= 3'b000;
      // memory_array[16196] <= 3'b000;
      // memory_array[16197] <= 3'b000;
      // memory_array[16198] <= 3'b110;
      // memory_array[16199] <= 3'b101;
      // memory_array[16200] <= 3'b000;
      // memory_array[16201] <= 3'b000;
      // memory_array[16202] <= 3'b000;
      // memory_array[16203] <= 3'b110;
      // memory_array[16204] <= 3'b110;
      // memory_array[16205] <= 3'b000;
      // memory_array[16206] <= 3'b000;
      // memory_array[16207] <= 3'b000;
      // memory_array[16208] <= 3'b101;
      // memory_array[16209] <= 3'b000;
      // memory_array[16210] <= 3'b000;
      // memory_array[16211] <= 3'b110;
      // memory_array[16212] <= 3'b111;
      // memory_array[16213] <= 3'b110;
      // memory_array[16214] <= 3'b110;
      // memory_array[16215] <= 3'b110;
      // memory_array[16216] <= 3'b111;
      // memory_array[16217] <= 3'b110;
      // memory_array[16218] <= 3'b110;
      // memory_array[16219] <= 3'b110;
      // memory_array[16220] <= 3'b110;
      // memory_array[16221] <= 3'b000;
      // memory_array[16222] <= 3'b000;
      // memory_array[16223] <= 3'b110;
      // memory_array[16224] <= 3'b110;
      // memory_array[16225] <= 3'b000;
      // memory_array[16226] <= 3'b111;
      // memory_array[16227] <= 3'b000;
      // memory_array[16228] <= 3'b110;
      // memory_array[16229] <= 3'b110;
      // memory_array[16230] <= 3'b110;
      // memory_array[16231] <= 3'b000;
      // memory_array[16232] <= 3'b000;
      // memory_array[16233] <= 3'b110;
      // memory_array[16234] <= 3'b110;
      // memory_array[16235] <= 3'b111;
      // memory_array[16236] <= 3'b111;
      // memory_array[16237] <= 3'b110;
      // memory_array[16238] <= 3'b000;
      // memory_array[16239] <= 3'b000;
      // memory_array[16240] <= 3'b111;
      // memory_array[16241] <= 3'b000;
      // memory_array[16242] <= 3'b000;
      // memory_array[16243] <= 3'b110;
      // memory_array[16244] <= 3'b111;
      // memory_array[16245] <= 3'b111;
      // memory_array[16246] <= 3'b111;
      // memory_array[16247] <= 3'b111;
      // memory_array[16248] <= 3'b111;
      // memory_array[16249] <= 3'b101;
      // memory_array[16250] <= 3'b000;
      // memory_array[16251] <= 3'b000;
      // memory_array[16252] <= 3'b000;
      // memory_array[16253] <= 3'b000;
      // memory_array[16254] <= 3'b111;
      // memory_array[16255] <= 3'b000;
      // memory_array[16256] <= 3'b000;
      // memory_array[16257] <= 3'b000;
      // memory_array[16258] <= 3'b000;
      // memory_array[16259] <= 3'b000;
      // memory_array[16260] <= 3'b111;
      // memory_array[16261] <= 3'b000;
      // memory_array[16262] <= 3'b000;
      // memory_array[16263] <= 3'b000;
      // memory_array[16264] <= 3'b000;
      // memory_array[16265] <= 3'b000;
      // memory_array[16266] <= 3'b000;
      // memory_array[16267] <= 3'b000;
      // memory_array[16268] <= 3'b000;
      // memory_array[16269] <= 3'b000;
      // memory_array[16270] <= 3'b000;
      // memory_array[16271] <= 3'b000;
      // memory_array[16272] <= 3'b000;
      // memory_array[16273] <= 3'b000;
      // memory_array[16274] <= 3'b000;
      // memory_array[16275] <= 3'b000;
      // memory_array[16276] <= 3'b000;
      // memory_array[16277] <= 3'b000;
      // memory_array[16278] <= 3'b000;
      // memory_array[16279] <= 3'b111;
      // memory_array[16280] <= 3'b000;
      // memory_array[16281] <= 3'b000;
      // memory_array[16282] <= 3'b000;
      // memory_array[16283] <= 3'b000;
      // memory_array[16284] <= 3'b000;
      // memory_array[16285] <= 3'b000;
      // memory_array[16286] <= 3'b000;
      // memory_array[16287] <= 3'b000;
      // memory_array[16288] <= 3'b110;
      // memory_array[16289] <= 3'b111;
      // memory_array[16290] <= 3'b111;
      // memory_array[16291] <= 3'b000;
      // memory_array[16292] <= 3'b000;
      // memory_array[16293] <= 3'b000;
      // memory_array[16294] <= 3'b000;
      // memory_array[16295] <= 3'b000;
      // memory_array[16296] <= 3'b000;
      // memory_array[16297] <= 3'b101;
      // memory_array[16298] <= 3'b101;
      // memory_array[16299] <= 3'b101;
      // memory_array[16300] <= 3'b000;
      // memory_array[16301] <= 3'b000;
      // memory_array[16302] <= 3'b000;
      // memory_array[16303] <= 3'b110;
      // memory_array[16304] <= 3'b101;
      // memory_array[16305] <= 3'b000;
      // memory_array[16306] <= 3'b000;
      // memory_array[16307] <= 3'b000;
      // memory_array[16308] <= 3'b000;
      // memory_array[16309] <= 3'b000;
      // memory_array[16310] <= 3'b000;
      // memory_array[16311] <= 3'b111;
      // memory_array[16312] <= 3'b000;
      // memory_array[16313] <= 3'b101;
      // memory_array[16314] <= 3'b000;
      // memory_array[16315] <= 3'b111;
      // memory_array[16316] <= 3'b000;
      // memory_array[16317] <= 3'b000;
      // memory_array[16318] <= 3'b000;
      // memory_array[16319] <= 3'b000;
      // memory_array[16320] <= 3'b000;
      // memory_array[16321] <= 3'b000;
      // memory_array[16322] <= 3'b000;
      // memory_array[16323] <= 3'b000;
      // memory_array[16324] <= 3'b000;
      // memory_array[16325] <= 3'b000;
      // memory_array[16326] <= 3'b000;
      // memory_array[16327] <= 3'b000;
      // memory_array[16328] <= 3'b000;
      // memory_array[16329] <= 3'b000;
      // memory_array[16330] <= 3'b000;
      // memory_array[16331] <= 3'b000;
      // memory_array[16332] <= 3'b000;
      // memory_array[16333] <= 3'b000;
      // memory_array[16334] <= 3'b000;
      // memory_array[16335] <= 3'b000;
      // memory_array[16336] <= 3'b000;
      // memory_array[16337] <= 3'b111;
      // memory_array[16338] <= 3'b111;
      // memory_array[16339] <= 3'b000;
      // memory_array[16340] <= 3'b000;
      // memory_array[16341] <= 3'b111;
      // memory_array[16342] <= 3'b000;
      // memory_array[16343] <= 3'b000;
      // memory_array[16344] <= 3'b000;
      // memory_array[16345] <= 3'b000;
      // memory_array[16346] <= 3'b000;
      // memory_array[16347] <= 3'b000;
      // memory_array[16348] <= 3'b000;
      // memory_array[16349] <= 3'b000;
      // memory_array[16350] <= 3'b111;
      // memory_array[16351] <= 3'b111;
      // memory_array[16352] <= 3'b000;
      // memory_array[16353] <= 3'b111;
      // memory_array[16354] <= 3'b000;
      // memory_array[16355] <= 3'b000;
      // memory_array[16356] <= 3'b110;
      // memory_array[16357] <= 3'b000;
      // memory_array[16358] <= 3'b110;
      // memory_array[16359] <= 3'b110;
      // memory_array[16360] <= 3'b000;
      // memory_array[16361] <= 3'b000;
      // memory_array[16362] <= 3'b110;
      // memory_array[16363] <= 3'b000;
      // memory_array[16364] <= 3'b111;
      // memory_array[16365] <= 3'b111;
      // memory_array[16366] <= 3'b110;
      // memory_array[16367] <= 3'b110;
      // memory_array[16368] <= 3'b110;
      // memory_array[16369] <= 3'b110;
      // memory_array[16370] <= 3'b000;
      // memory_array[16371] <= 3'b000;
      // memory_array[16372] <= 3'b000;
      // memory_array[16373] <= 3'b000;
      // memory_array[16374] <= 3'b111;
      // memory_array[16375] <= 3'b000;
      // memory_array[16376] <= 3'b110;
      // memory_array[16377] <= 3'b110;
      // memory_array[16378] <= 3'b000;
      // memory_array[16379] <= 3'b110;
      // memory_array[16380] <= 3'b111;
      // memory_array[16381] <= 3'b111;
      // memory_array[16382] <= 3'b111;
      // memory_array[16383] <= 3'b110;
      // memory_array[16384] <= 3'b110;
      // memory_array[16385] <= 3'b111;
      // memory_array[16386] <= 3'b111;
      // memory_array[16387] <= 3'b111;
      // memory_array[16388] <= 3'b110;
      // memory_array[16389] <= 3'b000;
      // memory_array[16390] <= 3'b000;
      // memory_array[16391] <= 3'b101;
      // memory_array[16392] <= 3'b000;
      // memory_array[16393] <= 3'b110;
      // memory_array[16394] <= 3'b110;
      // memory_array[16395] <= 3'b000;
      // memory_array[16396] <= 3'b000;
      // memory_array[16397] <= 3'b000;
      // memory_array[16398] <= 3'b110;
      // memory_array[16399] <= 3'b110;
      // memory_array[16400] <= 3'b101;
      // memory_array[16401] <= 3'b101;
      // memory_array[16402] <= 3'b101;
      // memory_array[16403] <= 3'b101;
      // memory_array[16404] <= 3'b101;
      // memory_array[16405] <= 3'b101;
      // memory_array[16406] <= 3'b101;
      // memory_array[16407] <= 3'b101;
      // memory_array[16408] <= 3'b101;
      // memory_array[16409] <= 3'b000;
      // memory_array[16410] <= 3'b000;
      // memory_array[16411] <= 3'b110;
      // memory_array[16412] <= 3'b111;
      // memory_array[16413] <= 3'b110;
      // memory_array[16414] <= 3'b110;
      // memory_array[16415] <= 3'b110;
      // memory_array[16416] <= 3'b111;
      // memory_array[16417] <= 3'b110;
      // memory_array[16418] <= 3'b110;
      // memory_array[16419] <= 3'b110;
      // memory_array[16420] <= 3'b110;
      // memory_array[16421] <= 3'b000;
      // memory_array[16422] <= 3'b000;
      // memory_array[16423] <= 3'b110;
      // memory_array[16424] <= 3'b000;
      // memory_array[16425] <= 3'b111;
      // memory_array[16426] <= 3'b111;
      // memory_array[16427] <= 3'b000;
      // memory_array[16428] <= 3'b110;
      // memory_array[16429] <= 3'b000;
      // memory_array[16430] <= 3'b111;
      // memory_array[16431] <= 3'b111;
      // memory_array[16432] <= 3'b111;
      // memory_array[16433] <= 3'b000;
      // memory_array[16434] <= 3'b110;
      // memory_array[16435] <= 3'b111;
      // memory_array[16436] <= 3'b000;
      // memory_array[16437] <= 3'b000;
      // memory_array[16438] <= 3'b111;
      // memory_array[16439] <= 3'b111;
      // memory_array[16440] <= 3'b111;
      // memory_array[16441] <= 3'b000;
      // memory_array[16442] <= 3'b000;
      // memory_array[16443] <= 3'b000;
      // memory_array[16444] <= 3'b111;
      // memory_array[16445] <= 3'b111;
      // memory_array[16446] <= 3'b000;
      // memory_array[16447] <= 3'b000;
      // memory_array[16448] <= 3'b000;
      // memory_array[16449] <= 3'b000;
      // memory_array[16450] <= 3'b000;
      // memory_array[16451] <= 3'b111;
      // memory_array[16452] <= 3'b111;
      // memory_array[16453] <= 3'b111;
      // memory_array[16454] <= 3'b111;
      // memory_array[16455] <= 3'b000;
      // memory_array[16456] <= 3'b000;
      // memory_array[16457] <= 3'b111;
      // memory_array[16458] <= 3'b111;
      // memory_array[16459] <= 3'b111;
      // memory_array[16460] <= 3'b111;
      // memory_array[16461] <= 3'b000;
      // memory_array[16462] <= 3'b000;
      // memory_array[16463] <= 3'b101;
      // memory_array[16464] <= 3'b111;
      // memory_array[16465] <= 3'b111;
      // memory_array[16466] <= 3'b111;
      // memory_array[16467] <= 3'b000;
      // memory_array[16468] <= 3'b000;
      // memory_array[16469] <= 3'b110;
      // memory_array[16470] <= 3'b000;
      // memory_array[16471] <= 3'b000;
      // memory_array[16472] <= 3'b000;
      // memory_array[16473] <= 3'b000;
      // memory_array[16474] <= 3'b000;
      // memory_array[16475] <= 3'b000;
      // memory_array[16476] <= 3'b000;
      // memory_array[16477] <= 3'b111;
      // memory_array[16478] <= 3'b111;
      // memory_array[16479] <= 3'b111;
      // memory_array[16480] <= 3'b111;
      // memory_array[16481] <= 3'b000;
      // memory_array[16482] <= 3'b000;
      // memory_array[16483] <= 3'b110;
      // memory_array[16484] <= 3'b000;
      // memory_array[16485] <= 3'b000;
      // memory_array[16486] <= 3'b000;
      // memory_array[16487] <= 3'b111;
      // memory_array[16488] <= 3'b111;
      // memory_array[16489] <= 3'b111;
      // memory_array[16490] <= 3'b111;
      // memory_array[16491] <= 3'b111;
      // memory_array[16492] <= 3'b000;
      // memory_array[16493] <= 3'b000;
      // memory_array[16494] <= 3'b000;
      // memory_array[16495] <= 3'b000;
      // memory_array[16496] <= 3'b000;
      // memory_array[16497] <= 3'b000;
      // memory_array[16498] <= 3'b000;
      // memory_array[16499] <= 3'b101;
      // memory_array[16500] <= 3'b000;
      // memory_array[16501] <= 3'b000;
      // memory_array[16502] <= 3'b000;
      // memory_array[16503] <= 3'b000;
      // memory_array[16504] <= 3'b110;
      // memory_array[16505] <= 3'b000;
      // memory_array[16506] <= 3'b000;
      // memory_array[16507] <= 3'b000;
      // memory_array[16508] <= 3'b000;
      // memory_array[16509] <= 3'b111;
      // memory_array[16510] <= 3'b111;
      // memory_array[16511] <= 3'b111;
      // memory_array[16512] <= 3'b111;
      // memory_array[16513] <= 3'b111;
      // memory_array[16514] <= 3'b111;
      // memory_array[16515] <= 3'b111;
      // memory_array[16516] <= 3'b111;
      // memory_array[16517] <= 3'b000;
      // memory_array[16518] <= 3'b000;
      // memory_array[16519] <= 3'b000;
      // memory_array[16520] <= 3'b000;
      // memory_array[16521] <= 3'b000;
      // memory_array[16522] <= 3'b000;
      // memory_array[16523] <= 3'b000;
      // memory_array[16524] <= 3'b101;
      // memory_array[16525] <= 3'b000;
      // memory_array[16526] <= 3'b111;
      // memory_array[16527] <= 3'b111;
      // memory_array[16528] <= 3'b111;
      // memory_array[16529] <= 3'b111;
      // memory_array[16530] <= 3'b111;
      // memory_array[16531] <= 3'b111;
      // memory_array[16532] <= 3'b000;
      // memory_array[16533] <= 3'b000;
      // memory_array[16534] <= 3'b000;
      // memory_array[16535] <= 3'b000;
      // memory_array[16536] <= 3'b111;
      // memory_array[16537] <= 3'b111;
      // memory_array[16538] <= 3'b111;
      // memory_array[16539] <= 3'b111;
      // memory_array[16540] <= 3'b111;
      // memory_array[16541] <= 3'b111;
      // memory_array[16542] <= 3'b111;
      // memory_array[16543] <= 3'b111;
      // memory_array[16544] <= 3'b000;
      // memory_array[16545] <= 3'b110;
      // memory_array[16546] <= 3'b110;
      // memory_array[16547] <= 3'b000;
      // memory_array[16548] <= 3'b101;
      // memory_array[16549] <= 3'b000;
      // memory_array[16550] <= 3'b000;
      // memory_array[16551] <= 3'b111;
      // memory_array[16552] <= 3'b111;
      // memory_array[16553] <= 3'b111;
      // memory_array[16554] <= 3'b111;
      // memory_array[16555] <= 3'b111;
      // memory_array[16556] <= 3'b111;
      // memory_array[16557] <= 3'b000;
      // memory_array[16558] <= 3'b110;
      // memory_array[16559] <= 3'b110;
      // memory_array[16560] <= 3'b000;
      // memory_array[16561] <= 3'b000;
      // memory_array[16562] <= 3'b111;
      // memory_array[16563] <= 3'b111;
      // memory_array[16564] <= 3'b111;
      // memory_array[16565] <= 3'b111;
      // memory_array[16566] <= 3'b000;
      // memory_array[16567] <= 3'b110;
      // memory_array[16568] <= 3'b110;
      // memory_array[16569] <= 3'b110;
      // memory_array[16570] <= 3'b000;
      // memory_array[16571] <= 3'b000;
      // memory_array[16572] <= 3'b111;
      // memory_array[16573] <= 3'b111;
      // memory_array[16574] <= 3'b111;
      // memory_array[16575] <= 3'b111;
      // memory_array[16576] <= 3'b000;
      // memory_array[16577] <= 3'b000;
      // memory_array[16578] <= 3'b000;
      // memory_array[16579] <= 3'b110;
      // memory_array[16580] <= 3'b111;
      // memory_array[16581] <= 3'b111;
      // memory_array[16582] <= 3'b111;
      // memory_array[16583] <= 3'b110;
      // memory_array[16584] <= 3'b110;
      // memory_array[16585] <= 3'b111;
      // memory_array[16586] <= 3'b111;
      // memory_array[16587] <= 3'b111;
      // memory_array[16588] <= 3'b110;
      // memory_array[16589] <= 3'b000;
      // memory_array[16590] <= 3'b000;
      // memory_array[16591] <= 3'b101;
      // memory_array[16592] <= 3'b101;
      // memory_array[16593] <= 3'b101;
      // memory_array[16594] <= 3'b101;
      // memory_array[16595] <= 3'b101;
      // memory_array[16596] <= 3'b101;
      // memory_array[16597] <= 3'b101;
      // memory_array[16598] <= 3'b101;
      // memory_array[16599] <= 3'b101;
      // memory_array[16600] <= 3'b101;
      // memory_array[16601] <= 3'b101;
      // memory_array[16602] <= 3'b101;
      // memory_array[16603] <= 3'b101;
      // memory_array[16604] <= 3'b101;
      // memory_array[16605] <= 3'b101;
      // memory_array[16606] <= 3'b101;
      // memory_array[16607] <= 3'b101;
      // memory_array[16608] <= 3'b101;
      // memory_array[16609] <= 3'b000;
      // memory_array[16610] <= 3'b000;
      // memory_array[16611] <= 3'b110;
      // memory_array[16612] <= 3'b110;
      // memory_array[16613] <= 3'b111;
      // memory_array[16614] <= 3'b111;
      // memory_array[16615] <= 3'b110;
      // memory_array[16616] <= 3'b110;
      // memory_array[16617] <= 3'b110;
      // memory_array[16618] <= 3'b110;
      // memory_array[16619] <= 3'b110;
      // memory_array[16620] <= 3'b110;
      // memory_array[16621] <= 3'b000;
      // memory_array[16622] <= 3'b000;
      // memory_array[16623] <= 3'b000;
      // memory_array[16624] <= 3'b111;
      // memory_array[16625] <= 3'b111;
      // memory_array[16626] <= 3'b111;
      // memory_array[16627] <= 3'b000;
      // memory_array[16628] <= 3'b000;
      // memory_array[16629] <= 3'b111;
      // memory_array[16630] <= 3'b111;
      // memory_array[16631] <= 3'b111;
      // memory_array[16632] <= 3'b111;
      // memory_array[16633] <= 3'b111;
      // memory_array[16634] <= 3'b111;
      // memory_array[16635] <= 3'b110;
      // memory_array[16636] <= 3'b000;
      // memory_array[16637] <= 3'b111;
      // memory_array[16638] <= 3'b111;
      // memory_array[16639] <= 3'b111;
      // memory_array[16640] <= 3'b111;
      // memory_array[16641] <= 3'b000;
      // memory_array[16642] <= 3'b000;
      // memory_array[16643] <= 3'b111;
      // memory_array[16644] <= 3'b111;
      // memory_array[16645] <= 3'b111;
      // memory_array[16646] <= 3'b000;
      // memory_array[16647] <= 3'b000;
      // memory_array[16648] <= 3'b000;
      // memory_array[16649] <= 3'b000;
      // memory_array[16650] <= 3'b111;
      // memory_array[16651] <= 3'b111;
      // memory_array[16652] <= 3'b111;
      // memory_array[16653] <= 3'b111;
      // memory_array[16654] <= 3'b111;
      // memory_array[16655] <= 3'b000;
      // memory_array[16656] <= 3'b111;
      // memory_array[16657] <= 3'b111;
      // memory_array[16658] <= 3'b111;
      // memory_array[16659] <= 3'b111;
      // memory_array[16660] <= 3'b111;
      // memory_array[16661] <= 3'b000;
      // memory_array[16662] <= 3'b000;
      // memory_array[16663] <= 3'b000;
      // memory_array[16664] <= 3'b111;
      // memory_array[16665] <= 3'b111;
      // memory_array[16666] <= 3'b111;
      // memory_array[16667] <= 3'b111;
      // memory_array[16668] <= 3'b111;
      // memory_array[16669] <= 3'b110;
      // memory_array[16670] <= 3'b000;
      // memory_array[16671] <= 3'b000;
      // memory_array[16672] <= 3'b000;
      // memory_array[16673] <= 3'b000;
      // memory_array[16674] <= 3'b000;
      // memory_array[16675] <= 3'b000;
      // memory_array[16676] <= 3'b111;
      // memory_array[16677] <= 3'b111;
      // memory_array[16678] <= 3'b111;
      // memory_array[16679] <= 3'b111;
      // memory_array[16680] <= 3'b111;
      // memory_array[16681] <= 3'b111;
      // memory_array[16682] <= 3'b000;
      // memory_array[16683] <= 3'b000;
      // memory_array[16684] <= 3'b000;
      // memory_array[16685] <= 3'b000;
      // memory_array[16686] <= 3'b000;
      // memory_array[16687] <= 3'b111;
      // memory_array[16688] <= 3'b111;
      // memory_array[16689] <= 3'b111;
      // memory_array[16690] <= 3'b111;
      // memory_array[16691] <= 3'b111;
      // memory_array[16692] <= 3'b111;
      // memory_array[16693] <= 3'b111;
      // memory_array[16694] <= 3'b000;
      // memory_array[16695] <= 3'b000;
      // memory_array[16696] <= 3'b000;
      // memory_array[16697] <= 3'b000;
      // memory_array[16698] <= 3'b000;
      // memory_array[16699] <= 3'b000;
      // memory_array[16700] <= 3'b000;
      // memory_array[16701] <= 3'b000;
      // memory_array[16702] <= 3'b110;
      // memory_array[16703] <= 3'b000;
      // memory_array[16704] <= 3'b000;
      // memory_array[16705] <= 3'b000;
      // memory_array[16706] <= 3'b000;
      // memory_array[16707] <= 3'b111;
      // memory_array[16708] <= 3'b111;
      // memory_array[16709] <= 3'b111;
      // memory_array[16710] <= 3'b111;
      // memory_array[16711] <= 3'b111;
      // memory_array[16712] <= 3'b111;
      // memory_array[16713] <= 3'b111;
      // memory_array[16714] <= 3'b111;
      // memory_array[16715] <= 3'b111;
      // memory_array[16716] <= 3'b111;
      // memory_array[16717] <= 3'b111;
      // memory_array[16718] <= 3'b000;
      // memory_array[16719] <= 3'b000;
      // memory_array[16720] <= 3'b000;
      // memory_array[16721] <= 3'b000;
      // memory_array[16722] <= 3'b000;
      // memory_array[16723] <= 3'b000;
      // memory_array[16724] <= 3'b000;
      // memory_array[16725] <= 3'b111;
      // memory_array[16726] <= 3'b111;
      // memory_array[16727] <= 3'b111;
      // memory_array[16728] <= 3'b111;
      // memory_array[16729] <= 3'b111;
      // memory_array[16730] <= 3'b111;
      // memory_array[16731] <= 3'b111;
      // memory_array[16732] <= 3'b111;
      // memory_array[16733] <= 3'b000;
      // memory_array[16734] <= 3'b111;
      // memory_array[16735] <= 3'b111;
      // memory_array[16736] <= 3'b111;
      // memory_array[16737] <= 3'b111;
      // memory_array[16738] <= 3'b111;
      // memory_array[16739] <= 3'b111;
      // memory_array[16740] <= 3'b111;
      // memory_array[16741] <= 3'b111;
      // memory_array[16742] <= 3'b111;
      // memory_array[16743] <= 3'b111;
      // memory_array[16744] <= 3'b111;
      // memory_array[16745] <= 3'b000;
      // memory_array[16746] <= 3'b101;
      // memory_array[16747] <= 3'b101;
      // memory_array[16748] <= 3'b000;
      // memory_array[16749] <= 3'b000;
      // memory_array[16750] <= 3'b111;
      // memory_array[16751] <= 3'b111;
      // memory_array[16752] <= 3'b111;
      // memory_array[16753] <= 3'b111;
      // memory_array[16754] <= 3'b111;
      // memory_array[16755] <= 3'b111;
      // memory_array[16756] <= 3'b111;
      // memory_array[16757] <= 3'b111;
      // memory_array[16758] <= 3'b000;
      // memory_array[16759] <= 3'b000;
      // memory_array[16760] <= 3'b000;
      // memory_array[16761] <= 3'b111;
      // memory_array[16762] <= 3'b111;
      // memory_array[16763] <= 3'b111;
      // memory_array[16764] <= 3'b111;
      // memory_array[16765] <= 3'b111;
      // memory_array[16766] <= 3'b110;
      // memory_array[16767] <= 3'b110;
      // memory_array[16768] <= 3'b000;
      // memory_array[16769] <= 3'b000;
      // memory_array[16770] <= 3'b110;
      // memory_array[16771] <= 3'b111;
      // memory_array[16772] <= 3'b111;
      // memory_array[16773] <= 3'b111;
      // memory_array[16774] <= 3'b111;
      // memory_array[16775] <= 3'b111;
      // memory_array[16776] <= 3'b111;
      // memory_array[16777] <= 3'b110;
      // memory_array[16778] <= 3'b000;
      // memory_array[16779] <= 3'b111;
      // memory_array[16780] <= 3'b110;
      // memory_array[16781] <= 3'b110;
      // memory_array[16782] <= 3'b110;
      // memory_array[16783] <= 3'b110;
      // memory_array[16784] <= 3'b110;
      // memory_array[16785] <= 3'b110;
      // memory_array[16786] <= 3'b110;
      // memory_array[16787] <= 3'b110;
      // memory_array[16788] <= 3'b110;
      // memory_array[16789] <= 3'b000;
      // memory_array[16790] <= 3'b000;
      // memory_array[16791] <= 3'b101;
      // memory_array[16792] <= 3'b101;
      // memory_array[16793] <= 3'b101;
      // memory_array[16794] <= 3'b101;
      // memory_array[16795] <= 3'b101;
      // memory_array[16796] <= 3'b101;
      // memory_array[16797] <= 3'b101;
      // memory_array[16798] <= 3'b101;
      // memory_array[16799] <= 3'b101;
      // memory_array[16800] <= 3'b000;
      // memory_array[16801] <= 3'b000;
      // memory_array[16802] <= 3'b000;
      // memory_array[16803] <= 3'b110;
      // memory_array[16804] <= 3'b110;
      // memory_array[16805] <= 3'b000;
      // memory_array[16806] <= 3'b000;
      // memory_array[16807] <= 3'b000;
      // memory_array[16808] <= 3'b101;
      // memory_array[16809] <= 3'b000;
      // memory_array[16810] <= 3'b000;
      // memory_array[16811] <= 3'b110;
      // memory_array[16812] <= 3'b111;
      // memory_array[16813] <= 3'b110;
      // memory_array[16814] <= 3'b110;
      // memory_array[16815] <= 3'b110;
      // memory_array[16816] <= 3'b111;
      // memory_array[16817] <= 3'b110;
      // memory_array[16818] <= 3'b110;
      // memory_array[16819] <= 3'b110;
      // memory_array[16820] <= 3'b000;
      // memory_array[16821] <= 3'b000;
      // memory_array[16822] <= 3'b111;
      // memory_array[16823] <= 3'b111;
      // memory_array[16824] <= 3'b111;
      // memory_array[16825] <= 3'b111;
      // memory_array[16826] <= 3'b111;
      // memory_array[16827] <= 3'b000;
      // memory_array[16828] <= 3'b111;
      // memory_array[16829] <= 3'b111;
      // memory_array[16830] <= 3'b111;
      // memory_array[16831] <= 3'b111;
      // memory_array[16832] <= 3'b111;
      // memory_array[16833] <= 3'b111;
      // memory_array[16834] <= 3'b000;
      // memory_array[16835] <= 3'b111;
      // memory_array[16836] <= 3'b000;
      // memory_array[16837] <= 3'b111;
      // memory_array[16838] <= 3'b111;
      // memory_array[16839] <= 3'b111;
      // memory_array[16840] <= 3'b111;
      // memory_array[16841] <= 3'b000;
      // memory_array[16842] <= 3'b111;
      // memory_array[16843] <= 3'b111;
      // memory_array[16844] <= 3'b111;
      // memory_array[16845] <= 3'b111;
      // memory_array[16846] <= 3'b111;
      // memory_array[16847] <= 3'b111;
      // memory_array[16848] <= 3'b110;
      // memory_array[16849] <= 3'b000;
      // memory_array[16850] <= 3'b000;
      // memory_array[16851] <= 3'b111;
      // memory_array[16852] <= 3'b111;
      // memory_array[16853] <= 3'b111;
      // memory_array[16854] <= 3'b111;
      // memory_array[16855] <= 3'b000;
      // memory_array[16856] <= 3'b000;
      // memory_array[16857] <= 3'b111;
      // memory_array[16858] <= 3'b111;
      // memory_array[16859] <= 3'b111;
      // memory_array[16860] <= 3'b111;
      // memory_array[16861] <= 3'b000;
      // memory_array[16862] <= 3'b111;
      // memory_array[16863] <= 3'b111;
      // memory_array[16864] <= 3'b111;
      // memory_array[16865] <= 3'b111;
      // memory_array[16866] <= 3'b111;
      // memory_array[16867] <= 3'b111;
      // memory_array[16868] <= 3'b111;
      // memory_array[16869] <= 3'b000;
      // memory_array[16870] <= 3'b000;
      // memory_array[16871] <= 3'b000;
      // memory_array[16872] <= 3'b000;
      // memory_array[16873] <= 3'b000;
      // memory_array[16874] <= 3'b000;
      // memory_array[16875] <= 3'b000;
      // memory_array[16876] <= 3'b111;
      // memory_array[16877] <= 3'b111;
      // memory_array[16878] <= 3'b111;
      // memory_array[16879] <= 3'b111;
      // memory_array[16880] <= 3'b111;
      // memory_array[16881] <= 3'b111;
      // memory_array[16882] <= 3'b111;
      // memory_array[16883] <= 3'b000;
      // memory_array[16884] <= 3'b000;
      // memory_array[16885] <= 3'b000;
      // memory_array[16886] <= 3'b111;
      // memory_array[16887] <= 3'b111;
      // memory_array[16888] <= 3'b111;
      // memory_array[16889] <= 3'b111;
      // memory_array[16890] <= 3'b111;
      // memory_array[16891] <= 3'b111;
      // memory_array[16892] <= 3'b111;
      // memory_array[16893] <= 3'b111;
      // memory_array[16894] <= 3'b000;
      // memory_array[16895] <= 3'b000;
      // memory_array[16896] <= 3'b000;
      // memory_array[16897] <= 3'b000;
      // memory_array[16898] <= 3'b000;
      // memory_array[16899] <= 3'b000;
      // memory_array[16900] <= 3'b000;
      // memory_array[16901] <= 3'b000;
      // memory_array[16902] <= 3'b000;
      // memory_array[16903] <= 3'b000;
      // memory_array[16904] <= 3'b000;
      // memory_array[16905] <= 3'b000;
      // memory_array[16906] <= 3'b111;
      // memory_array[16907] <= 3'b111;
      // memory_array[16908] <= 3'b111;
      // memory_array[16909] <= 3'b111;
      // memory_array[16910] <= 3'b111;
      // memory_array[16911] <= 3'b111;
      // memory_array[16912] <= 3'b111;
      // memory_array[16913] <= 3'b111;
      // memory_array[16914] <= 3'b000;
      // memory_array[16915] <= 3'b111;
      // memory_array[16916] <= 3'b111;
      // memory_array[16917] <= 3'b111;
      // memory_array[16918] <= 3'b111;
      // memory_array[16919] <= 3'b000;
      // memory_array[16920] <= 3'b000;
      // memory_array[16921] <= 3'b000;
      // memory_array[16922] <= 3'b000;
      // memory_array[16923] <= 3'b000;
      // memory_array[16924] <= 3'b111;
      // memory_array[16925] <= 3'b111;
      // memory_array[16926] <= 3'b111;
      // memory_array[16927] <= 3'b111;
      // memory_array[16928] <= 3'b111;
      // memory_array[16929] <= 3'b111;
      // memory_array[16930] <= 3'b111;
      // memory_array[16931] <= 3'b111;
      // memory_array[16932] <= 3'b111;
      // memory_array[16933] <= 3'b111;
      // memory_array[16934] <= 3'b000;
      // memory_array[16935] <= 3'b111;
      // memory_array[16936] <= 3'b111;
      // memory_array[16937] <= 3'b111;
      // memory_array[16938] <= 3'b111;
      // memory_array[16939] <= 3'b111;
      // memory_array[16940] <= 3'b111;
      // memory_array[16941] <= 3'b111;
      // memory_array[16942] <= 3'b111;
      // memory_array[16943] <= 3'b111;
      // memory_array[16944] <= 3'b111;
      // memory_array[16945] <= 3'b111;
      // memory_array[16946] <= 3'b110;
      // memory_array[16947] <= 3'b110;
      // memory_array[16948] <= 3'b101;
      // memory_array[16949] <= 3'b111;
      // memory_array[16950] <= 3'b111;
      // memory_array[16951] <= 3'b111;
      // memory_array[16952] <= 3'b111;
      // memory_array[16953] <= 3'b111;
      // memory_array[16954] <= 3'b111;
      // memory_array[16955] <= 3'b111;
      // memory_array[16956] <= 3'b111;
      // memory_array[16957] <= 3'b111;
      // memory_array[16958] <= 3'b111;
      // memory_array[16959] <= 3'b000;
      // memory_array[16960] <= 3'b000;
      // memory_array[16961] <= 3'b111;
      // memory_array[16962] <= 3'b111;
      // memory_array[16963] <= 3'b111;
      // memory_array[16964] <= 3'b111;
      // memory_array[16965] <= 3'b111;
      // memory_array[16966] <= 3'b000;
      // memory_array[16967] <= 3'b110;
      // memory_array[16968] <= 3'b110;
      // memory_array[16969] <= 3'b110;
      // memory_array[16970] <= 3'b000;
      // memory_array[16971] <= 3'b111;
      // memory_array[16972] <= 3'b111;
      // memory_array[16973] <= 3'b111;
      // memory_array[16974] <= 3'b111;
      // memory_array[16975] <= 3'b111;
      // memory_array[16976] <= 3'b111;
      // memory_array[16977] <= 3'b000;
      // memory_array[16978] <= 3'b000;
      // memory_array[16979] <= 3'b110;
      // memory_array[16980] <= 3'b111;
      // memory_array[16981] <= 3'b111;
      // memory_array[16982] <= 3'b111;
      // memory_array[16983] <= 3'b110;
      // memory_array[16984] <= 3'b110;
      // memory_array[16985] <= 3'b111;
      // memory_array[16986] <= 3'b111;
      // memory_array[16987] <= 3'b111;
      // memory_array[16988] <= 3'b110;
      // memory_array[16989] <= 3'b000;
      // memory_array[16990] <= 3'b000;
      // memory_array[16991] <= 3'b101;
      // memory_array[16992] <= 3'b000;
      // memory_array[16993] <= 3'b110;
      // memory_array[16994] <= 3'b110;
      // memory_array[16995] <= 3'b000;
      // memory_array[16996] <= 3'b000;
      // memory_array[16997] <= 3'b000;
      // memory_array[16998] <= 3'b110;
      // memory_array[16999] <= 3'b110;
      // memory_array[17000] <= 3'b101;
      // memory_array[17001] <= 3'b110;
      // memory_array[17002] <= 3'b110;
      // memory_array[17003] <= 3'b000;
      // memory_array[17004] <= 3'b000;
      // memory_array[17005] <= 3'b110;
      // memory_array[17006] <= 3'b110;
      // memory_array[17007] <= 3'b101;
      // memory_array[17008] <= 3'b101;
      // memory_array[17009] <= 3'b000;
      // memory_array[17010] <= 3'b000;
      // memory_array[17011] <= 3'b110;
      // memory_array[17012] <= 3'b110;
      // memory_array[17013] <= 3'b110;
      // memory_array[17014] <= 3'b110;
      // memory_array[17015] <= 3'b110;
      // memory_array[17016] <= 3'b110;
      // memory_array[17017] <= 3'b110;
      // memory_array[17018] <= 3'b000;
      // memory_array[17019] <= 3'b000;
      // memory_array[17020] <= 3'b000;
      // memory_array[17021] <= 3'b111;
      // memory_array[17022] <= 3'b111;
      // memory_array[17023] <= 3'b111;
      // memory_array[17024] <= 3'b111;
      // memory_array[17025] <= 3'b111;
      // memory_array[17026] <= 3'b111;
      // memory_array[17027] <= 3'b111;
      // memory_array[17028] <= 3'b111;
      // memory_array[17029] <= 3'b111;
      // memory_array[17030] <= 3'b111;
      // memory_array[17031] <= 3'b111;
      // memory_array[17032] <= 3'b111;
      // memory_array[17033] <= 3'b111;
      // memory_array[17034] <= 3'b111;
      // memory_array[17035] <= 3'b000;
      // memory_array[17036] <= 3'b110;
      // memory_array[17037] <= 3'b111;
      // memory_array[17038] <= 3'b111;
      // memory_array[17039] <= 3'b111;
      // memory_array[17040] <= 3'b111;
      // memory_array[17041] <= 3'b111;
      // memory_array[17042] <= 3'b111;
      // memory_array[17043] <= 3'b111;
      // memory_array[17044] <= 3'b111;
      // memory_array[17045] <= 3'b111;
      // memory_array[17046] <= 3'b111;
      // memory_array[17047] <= 3'b000;
      // memory_array[17048] <= 3'b000;
      // memory_array[17049] <= 3'b000;
      // memory_array[17050] <= 3'b000;
      // memory_array[17051] <= 3'b111;
      // memory_array[17052] <= 3'b111;
      // memory_array[17053] <= 3'b111;
      // memory_array[17054] <= 3'b111;
      // memory_array[17055] <= 3'b000;
      // memory_array[17056] <= 3'b000;
      // memory_array[17057] <= 3'b111;
      // memory_array[17058] <= 3'b111;
      // memory_array[17059] <= 3'b111;
      // memory_array[17060] <= 3'b111;
      // memory_array[17061] <= 3'b111;
      // memory_array[17062] <= 3'b111;
      // memory_array[17063] <= 3'b111;
      // memory_array[17064] <= 3'b111;
      // memory_array[17065] <= 3'b111;
      // memory_array[17066] <= 3'b111;
      // memory_array[17067] <= 3'b111;
      // memory_array[17068] <= 3'b111;
      // memory_array[17069] <= 3'b111;
      // memory_array[17070] <= 3'b000;
      // memory_array[17071] <= 3'b000;
      // memory_array[17072] <= 3'b000;
      // memory_array[17073] <= 3'b000;
      // memory_array[17074] <= 3'b111;
      // memory_array[17075] <= 3'b111;
      // memory_array[17076] <= 3'b111;
      // memory_array[17077] <= 3'b111;
      // memory_array[17078] <= 3'b000;
      // memory_array[17079] <= 3'b111;
      // memory_array[17080] <= 3'b111;
      // memory_array[17081] <= 3'b111;
      // memory_array[17082] <= 3'b111;
      // memory_array[17083] <= 3'b111;
      // memory_array[17084] <= 3'b000;
      // memory_array[17085] <= 3'b111;
      // memory_array[17086] <= 3'b111;
      // memory_array[17087] <= 3'b111;
      // memory_array[17088] <= 3'b111;
      // memory_array[17089] <= 3'b000;
      // memory_array[17090] <= 3'b111;
      // memory_array[17091] <= 3'b111;
      // memory_array[17092] <= 3'b111;
      // memory_array[17093] <= 3'b111;
      // memory_array[17094] <= 3'b111;
      // memory_array[17095] <= 3'b000;
      // memory_array[17096] <= 3'b000;
      // memory_array[17097] <= 3'b000;
      // memory_array[17098] <= 3'b000;
      // memory_array[17099] <= 3'b000;
      // memory_array[17100] <= 3'b000;
      // memory_array[17101] <= 3'b000;
      // memory_array[17102] <= 3'b000;
      // memory_array[17103] <= 3'b000;
      // memory_array[17104] <= 3'b000;
      // memory_array[17105] <= 3'b000;
      // memory_array[17106] <= 3'b000;
      // memory_array[17107] <= 3'b111;
      // memory_array[17108] <= 3'b111;
      // memory_array[17109] <= 3'b111;
      // memory_array[17110] <= 3'b111;
      // memory_array[17111] <= 3'b111;
      // memory_array[17112] <= 3'b111;
      // memory_array[17113] <= 3'b000;
      // memory_array[17114] <= 3'b000;
      // memory_array[17115] <= 3'b000;
      // memory_array[17116] <= 3'b111;
      // memory_array[17117] <= 3'b111;
      // memory_array[17118] <= 3'b111;
      // memory_array[17119] <= 3'b000;
      // memory_array[17120] <= 3'b000;
      // memory_array[17121] <= 3'b000;
      // memory_array[17122] <= 3'b111;
      // memory_array[17123] <= 3'b111;
      // memory_array[17124] <= 3'b111;
      // memory_array[17125] <= 3'b111;
      // memory_array[17126] <= 3'b111;
      // memory_array[17127] <= 3'b000;
      // memory_array[17128] <= 3'b111;
      // memory_array[17129] <= 3'b111;
      // memory_array[17130] <= 3'b111;
      // memory_array[17131] <= 3'b111;
      // memory_array[17132] <= 3'b111;
      // memory_array[17133] <= 3'b000;
      // memory_array[17134] <= 3'b000;
      // memory_array[17135] <= 3'b111;
      // memory_array[17136] <= 3'b111;
      // memory_array[17137] <= 3'b111;
      // memory_array[17138] <= 3'b111;
      // memory_array[17139] <= 3'b111;
      // memory_array[17140] <= 3'b000;
      // memory_array[17141] <= 3'b111;
      // memory_array[17142] <= 3'b111;
      // memory_array[17143] <= 3'b111;
      // memory_array[17144] <= 3'b111;
      // memory_array[17145] <= 3'b111;
      // memory_array[17146] <= 3'b000;
      // memory_array[17147] <= 3'b101;
      // memory_array[17148] <= 3'b000;
      // memory_array[17149] <= 3'b111;
      // memory_array[17150] <= 3'b111;
      // memory_array[17151] <= 3'b111;
      // memory_array[17152] <= 3'b000;
      // memory_array[17153] <= 3'b111;
      // memory_array[17154] <= 3'b111;
      // memory_array[17155] <= 3'b111;
      // memory_array[17156] <= 3'b111;
      // memory_array[17157] <= 3'b111;
      // memory_array[17158] <= 3'b111;
      // memory_array[17159] <= 3'b111;
      // memory_array[17160] <= 3'b000;
      // memory_array[17161] <= 3'b000;
      // memory_array[17162] <= 3'b111;
      // memory_array[17163] <= 3'b111;
      // memory_array[17164] <= 3'b111;
      // memory_array[17165] <= 3'b111;
      // memory_array[17166] <= 3'b000;
      // memory_array[17167] <= 3'b110;
      // memory_array[17168] <= 3'b000;
      // memory_array[17169] <= 3'b000;
      // memory_array[17170] <= 3'b111;
      // memory_array[17171] <= 3'b111;
      // memory_array[17172] <= 3'b111;
      // memory_array[17173] <= 3'b111;
      // memory_array[17174] <= 3'b111;
      // memory_array[17175] <= 3'b111;
      // memory_array[17176] <= 3'b111;
      // memory_array[17177] <= 3'b111;
      // memory_array[17178] <= 3'b000;
      // memory_array[17179] <= 3'b111;
      // memory_array[17180] <= 3'b110;
      // memory_array[17181] <= 3'b110;
      // memory_array[17182] <= 3'b110;
      // memory_array[17183] <= 3'b000;
      // memory_array[17184] <= 3'b111;
      // memory_array[17185] <= 3'b110;
      // memory_array[17186] <= 3'b110;
      // memory_array[17187] <= 3'b110;
      // memory_array[17188] <= 3'b000;
      // memory_array[17189] <= 3'b000;
      // memory_array[17190] <= 3'b000;
      // memory_array[17191] <= 3'b101;
      // memory_array[17192] <= 3'b110;
      // memory_array[17193] <= 3'b000;
      // memory_array[17194] <= 3'b000;
      // memory_array[17195] <= 3'b110;
      // memory_array[17196] <= 3'b110;
      // memory_array[17197] <= 3'b110;
      // memory_array[17198] <= 3'b000;
      // memory_array[17199] <= 3'b101;
      // memory_array[17200] <= 3'b101;
      // memory_array[17201] <= 3'b101;
      // memory_array[17202] <= 3'b110;
      // memory_array[17203] <= 3'b101;
      // memory_array[17204] <= 3'b101;
      // memory_array[17205] <= 3'b110;
      // memory_array[17206] <= 3'b101;
      // memory_array[17207] <= 3'b101;
      // memory_array[17208] <= 3'b101;
      // memory_array[17209] <= 3'b000;
      // memory_array[17210] <= 3'b000;
      // memory_array[17211] <= 3'b110;
      // memory_array[17212] <= 3'b110;
      // memory_array[17213] <= 3'b110;
      // memory_array[17214] <= 3'b110;
      // memory_array[17215] <= 3'b110;
      // memory_array[17216] <= 3'b110;
      // memory_array[17217] <= 3'b110;
      // memory_array[17218] <= 3'b110;
      // memory_array[17219] <= 3'b110;
      // memory_array[17220] <= 3'b110;
      // memory_array[17221] <= 3'b000;
      // memory_array[17222] <= 3'b000;
      // memory_array[17223] <= 3'b000;
      // memory_array[17224] <= 3'b111;
      // memory_array[17225] <= 3'b111;
      // memory_array[17226] <= 3'b111;
      // memory_array[17227] <= 3'b111;
      // memory_array[17228] <= 3'b111;
      // memory_array[17229] <= 3'b110;
      // memory_array[17230] <= 3'b110;
      // memory_array[17231] <= 3'b000;
      // memory_array[17232] <= 3'b111;
      // memory_array[17233] <= 3'b111;
      // memory_array[17234] <= 3'b111;
      // memory_array[17235] <= 3'b111;
      // memory_array[17236] <= 3'b110;
      // memory_array[17237] <= 3'b111;
      // memory_array[17238] <= 3'b111;
      // memory_array[17239] <= 3'b111;
      // memory_array[17240] <= 3'b111;
      // memory_array[17241] <= 3'b111;
      // memory_array[17242] <= 3'b000;
      // memory_array[17243] <= 3'b000;
      // memory_array[17244] <= 3'b111;
      // memory_array[17245] <= 3'b111;
      // memory_array[17246] <= 3'b111;
      // memory_array[17247] <= 3'b111;
      // memory_array[17248] <= 3'b000;
      // memory_array[17249] <= 3'b000;
      // memory_array[17250] <= 3'b000;
      // memory_array[17251] <= 3'b111;
      // memory_array[17252] <= 3'b111;
      // memory_array[17253] <= 3'b111;
      // memory_array[17254] <= 3'b111;
      // memory_array[17255] <= 3'b000;
      // memory_array[17256] <= 3'b110;
      // memory_array[17257] <= 3'b111;
      // memory_array[17258] <= 3'b111;
      // memory_array[17259] <= 3'b111;
      // memory_array[17260] <= 3'b111;
      // memory_array[17261] <= 3'b111;
      // memory_array[17262] <= 3'b000;
      // memory_array[17263] <= 3'b000;
      // memory_array[17264] <= 3'b000;
      // memory_array[17265] <= 3'b000;
      // memory_array[17266] <= 3'b111;
      // memory_array[17267] <= 3'b111;
      // memory_array[17268] <= 3'b111;
      // memory_array[17269] <= 3'b111;
      // memory_array[17270] <= 3'b111;
      // memory_array[17271] <= 3'b000;
      // memory_array[17272] <= 3'b000;
      // memory_array[17273] <= 3'b111;
      // memory_array[17274] <= 3'b111;
      // memory_array[17275] <= 3'b111;
      // memory_array[17276] <= 3'b111;
      // memory_array[17277] <= 3'b000;
      // memory_array[17278] <= 3'b000;
      // memory_array[17279] <= 3'b000;
      // memory_array[17280] <= 3'b110;
      // memory_array[17281] <= 3'b111;
      // memory_array[17282] <= 3'b111;
      // memory_array[17283] <= 3'b000;
      // memory_array[17284] <= 3'b111;
      // memory_array[17285] <= 3'b111;
      // memory_array[17286] <= 3'b111;
      // memory_array[17287] <= 3'b000;
      // memory_array[17288] <= 3'b000;
      // memory_array[17289] <= 3'b000;
      // memory_array[17290] <= 3'b000;
      // memory_array[17291] <= 3'b000;
      // memory_array[17292] <= 3'b111;
      // memory_array[17293] <= 3'b111;
      // memory_array[17294] <= 3'b000;
      // memory_array[17295] <= 3'b000;
      // memory_array[17296] <= 3'b000;
      // memory_array[17297] <= 3'b101;
      // memory_array[17298] <= 3'b000;
      // memory_array[17299] <= 3'b000;
      // memory_array[17300] <= 3'b101;
      // memory_array[17301] <= 3'b000;
      // memory_array[17302] <= 3'b000;
      // memory_array[17303] <= 3'b111;
      // memory_array[17304] <= 3'b111;
      // memory_array[17305] <= 3'b111;
      // memory_array[17306] <= 3'b111;
      // memory_array[17307] <= 3'b000;
      // memory_array[17308] <= 3'b111;
      // memory_array[17309] <= 3'b111;
      // memory_array[17310] <= 3'b111;
      // memory_array[17311] <= 3'b111;
      // memory_array[17312] <= 3'b000;
      // memory_array[17313] <= 3'b000;
      // memory_array[17314] <= 3'b000;
      // memory_array[17315] <= 3'b000;
      // memory_array[17316] <= 3'b111;
      // memory_array[17317] <= 3'b111;
      // memory_array[17318] <= 3'b111;
      // memory_array[17319] <= 3'b111;
      // memory_array[17320] <= 3'b000;
      // memory_array[17321] <= 3'b000;
      // memory_array[17322] <= 3'b111;
      // memory_array[17323] <= 3'b111;
      // memory_array[17324] <= 3'b111;
      // memory_array[17325] <= 3'b111;
      // memory_array[17326] <= 3'b000;
      // memory_array[17327] <= 3'b000;
      // memory_array[17328] <= 3'b000;
      // memory_array[17329] <= 3'b000;
      // memory_array[17330] <= 3'b000;
      // memory_array[17331] <= 3'b111;
      // memory_array[17332] <= 3'b000;
      // memory_array[17333] <= 3'b000;
      // memory_array[17334] <= 3'b000;
      // memory_array[17335] <= 3'b111;
      // memory_array[17336] <= 3'b111;
      // memory_array[17337] <= 3'b111;
      // memory_array[17338] <= 3'b111;
      // memory_array[17339] <= 3'b000;
      // memory_array[17340] <= 3'b101;
      // memory_array[17341] <= 3'b101;
      // memory_array[17342] <= 3'b111;
      // memory_array[17343] <= 3'b111;
      // memory_array[17344] <= 3'b111;
      // memory_array[17345] <= 3'b111;
      // memory_array[17346] <= 3'b111;
      // memory_array[17347] <= 3'b000;
      // memory_array[17348] <= 3'b111;
      // memory_array[17349] <= 3'b111;
      // memory_array[17350] <= 3'b111;
      // memory_array[17351] <= 3'b111;
      // memory_array[17352] <= 3'b000;
      // memory_array[17353] <= 3'b000;
      // memory_array[17354] <= 3'b000;
      // memory_array[17355] <= 3'b000;
      // memory_array[17356] <= 3'b111;
      // memory_array[17357] <= 3'b111;
      // memory_array[17358] <= 3'b111;
      // memory_array[17359] <= 3'b000;
      // memory_array[17360] <= 3'b110;
      // memory_array[17361] <= 3'b000;
      // memory_array[17362] <= 3'b111;
      // memory_array[17363] <= 3'b111;
      // memory_array[17364] <= 3'b111;
      // memory_array[17365] <= 3'b111;
      // memory_array[17366] <= 3'b110;
      // memory_array[17367] <= 3'b110;
      // memory_array[17368] <= 3'b000;
      // memory_array[17369] <= 3'b111;
      // memory_array[17370] <= 3'b111;
      // memory_array[17371] <= 3'b111;
      // memory_array[17372] <= 3'b000;
      // memory_array[17373] <= 3'b111;
      // memory_array[17374] <= 3'b111;
      // memory_array[17375] <= 3'b111;
      // memory_array[17376] <= 3'b111;
      // memory_array[17377] <= 3'b111;
      // memory_array[17378] <= 3'b111;
      // memory_array[17379] <= 3'b111;
      // memory_array[17380] <= 3'b110;
      // memory_array[17381] <= 3'b110;
      // memory_array[17382] <= 3'b110;
      // memory_array[17383] <= 3'b110;
      // memory_array[17384] <= 3'b111;
      // memory_array[17385] <= 3'b110;
      // memory_array[17386] <= 3'b110;
      // memory_array[17387] <= 3'b110;
      // memory_array[17388] <= 3'b111;
      // memory_array[17389] <= 3'b000;
      // memory_array[17390] <= 3'b000;
      // memory_array[17391] <= 3'b101;
      // memory_array[17392] <= 3'b101;
      // memory_array[17393] <= 3'b101;
      // memory_array[17394] <= 3'b000;
      // memory_array[17395] <= 3'b101;
      // memory_array[17396] <= 3'b101;
      // memory_array[17397] <= 3'b110;
      // memory_array[17398] <= 3'b101;
      // memory_array[17399] <= 3'b101;
      // memory_array[17400] <= 3'b101;
      // memory_array[17401] <= 3'b101;
      // memory_array[17402] <= 3'b101;
      // memory_array[17403] <= 3'b111;
      // memory_array[17404] <= 3'b111;
      // memory_array[17405] <= 3'b101;
      // memory_array[17406] <= 3'b101;
      // memory_array[17407] <= 3'b101;
      // memory_array[17408] <= 3'b101;
      // memory_array[17409] <= 3'b000;
      // memory_array[17410] <= 3'b000;
      // memory_array[17411] <= 3'b110;
      // memory_array[17412] <= 3'b111;
      // memory_array[17413] <= 3'b110;
      // memory_array[17414] <= 3'b110;
      // memory_array[17415] <= 3'b110;
      // memory_array[17416] <= 3'b110;
      // memory_array[17417] <= 3'b111;
      // memory_array[17418] <= 3'b110;
      // memory_array[17419] <= 3'b110;
      // memory_array[17420] <= 3'b111;
      // memory_array[17421] <= 3'b000;
      // memory_array[17422] <= 3'b110;
      // memory_array[17423] <= 3'b000;
      // memory_array[17424] <= 3'b111;
      // memory_array[17425] <= 3'b111;
      // memory_array[17426] <= 3'b111;
      // memory_array[17427] <= 3'b111;
      // memory_array[17428] <= 3'b000;
      // memory_array[17429] <= 3'b110;
      // memory_array[17430] <= 3'b111;
      // memory_array[17431] <= 3'b111;
      // memory_array[17432] <= 3'b111;
      // memory_array[17433] <= 3'b111;
      // memory_array[17434] <= 3'b111;
      // memory_array[17435] <= 3'b111;
      // memory_array[17436] <= 3'b110;
      // memory_array[17437] <= 3'b111;
      // memory_array[17438] <= 3'b111;
      // memory_array[17439] <= 3'b111;
      // memory_array[17440] <= 3'b111;
      // memory_array[17441] <= 3'b111;
      // memory_array[17442] <= 3'b000;
      // memory_array[17443] <= 3'b000;
      // memory_array[17444] <= 3'b000;
      // memory_array[17445] <= 3'b111;
      // memory_array[17446] <= 3'b111;
      // memory_array[17447] <= 3'b111;
      // memory_array[17448] <= 3'b111;
      // memory_array[17449] <= 3'b000;
      // memory_array[17450] <= 3'b000;
      // memory_array[17451] <= 3'b111;
      // memory_array[17452] <= 3'b111;
      // memory_array[17453] <= 3'b111;
      // memory_array[17454] <= 3'b111;
      // memory_array[17455] <= 3'b000;
      // memory_array[17456] <= 3'b000;
      // memory_array[17457] <= 3'b111;
      // memory_array[17458] <= 3'b111;
      // memory_array[17459] <= 3'b111;
      // memory_array[17460] <= 3'b111;
      // memory_array[17461] <= 3'b111;
      // memory_array[17462] <= 3'b000;
      // memory_array[17463] <= 3'b101;
      // memory_array[17464] <= 3'b101;
      // memory_array[17465] <= 3'b000;
      // memory_array[17466] <= 3'b000;
      // memory_array[17467] <= 3'b111;
      // memory_array[17468] <= 3'b111;
      // memory_array[17469] <= 3'b111;
      // memory_array[17470] <= 3'b111;
      // memory_array[17471] <= 3'b000;
      // memory_array[17472] <= 3'b000;
      // memory_array[17473] <= 3'b111;
      // memory_array[17474] <= 3'b111;
      // memory_array[17475] <= 3'b111;
      // memory_array[17476] <= 3'b000;
      // memory_array[17477] <= 3'b000;
      // memory_array[17478] <= 3'b000;
      // memory_array[17479] <= 3'b101;
      // memory_array[17480] <= 3'b000;
      // memory_array[17481] <= 3'b000;
      // memory_array[17482] <= 3'b000;
      // memory_array[17483] <= 3'b000;
      // memory_array[17484] <= 3'b111;
      // memory_array[17485] <= 3'b111;
      // memory_array[17486] <= 3'b111;
      // memory_array[17487] <= 3'b000;
      // memory_array[17488] <= 3'b000;
      // memory_array[17489] <= 3'b000;
      // memory_array[17490] <= 3'b000;
      // memory_array[17491] <= 3'b000;
      // memory_array[17492] <= 3'b000;
      // memory_array[17493] <= 3'b111;
      // memory_array[17494] <= 3'b000;
      // memory_array[17495] <= 3'b000;
      // memory_array[17496] <= 3'b000;
      // memory_array[17497] <= 3'b110;
      // memory_array[17498] <= 3'b110;
      // memory_array[17499] <= 3'b110;
      // memory_array[17500] <= 3'b000;
      // memory_array[17501] <= 3'b000;
      // memory_array[17502] <= 3'b111;
      // memory_array[17503] <= 3'b111;
      // memory_array[17504] <= 3'b000;
      // memory_array[17505] <= 3'b000;
      // memory_array[17506] <= 3'b111;
      // memory_array[17507] <= 3'b000;
      // memory_array[17508] <= 3'b111;
      // memory_array[17509] <= 3'b111;
      // memory_array[17510] <= 3'b111;
      // memory_array[17511] <= 3'b111;
      // memory_array[17512] <= 3'b000;
      // memory_array[17513] <= 3'b000;
      // memory_array[17514] <= 3'b000;
      // memory_array[17515] <= 3'b000;
      // memory_array[17516] <= 3'b000;
      // memory_array[17517] <= 3'b111;
      // memory_array[17518] <= 3'b111;
      // memory_array[17519] <= 3'b111;
      // memory_array[17520] <= 3'b000;
      // memory_array[17521] <= 3'b000;
      // memory_array[17522] <= 3'b111;
      // memory_array[17523] <= 3'b111;
      // memory_array[17524] <= 3'b111;
      // memory_array[17525] <= 3'b111;
      // memory_array[17526] <= 3'b000;
      // memory_array[17527] <= 3'b000;
      // memory_array[17528] <= 3'b000;
      // memory_array[17529] <= 3'b000;
      // memory_array[17530] <= 3'b000;
      // memory_array[17531] <= 3'b111;
      // memory_array[17532] <= 3'b000;
      // memory_array[17533] <= 3'b110;
      // memory_array[17534] <= 3'b000;
      // memory_array[17535] <= 3'b111;
      // memory_array[17536] <= 3'b111;
      // memory_array[17537] <= 3'b111;
      // memory_array[17538] <= 3'b111;
      // memory_array[17539] <= 3'b000;
      // memory_array[17540] <= 3'b000;
      // memory_array[17541] <= 3'b000;
      // memory_array[17542] <= 3'b111;
      // memory_array[17543] <= 3'b111;
      // memory_array[17544] <= 3'b111;
      // memory_array[17545] <= 3'b111;
      // memory_array[17546] <= 3'b111;
      // memory_array[17547] <= 3'b000;
      // memory_array[17548] <= 3'b111;
      // memory_array[17549] <= 3'b111;
      // memory_array[17550] <= 3'b111;
      // memory_array[17551] <= 3'b111;
      // memory_array[17552] <= 3'b000;
      // memory_array[17553] <= 3'b000;
      // memory_array[17554] <= 3'b110;
      // memory_array[17555] <= 3'b000;
      // memory_array[17556] <= 3'b000;
      // memory_array[17557] <= 3'b111;
      // memory_array[17558] <= 3'b000;
      // memory_array[17559] <= 3'b000;
      // memory_array[17560] <= 3'b000;
      // memory_array[17561] <= 3'b000;
      // memory_array[17562] <= 3'b111;
      // memory_array[17563] <= 3'b111;
      // memory_array[17564] <= 3'b111;
      // memory_array[17565] <= 3'b111;
      // memory_array[17566] <= 3'b110;
      // memory_array[17567] <= 3'b000;
      // memory_array[17568] <= 3'b111;
      // memory_array[17569] <= 3'b111;
      // memory_array[17570] <= 3'b111;
      // memory_array[17571] <= 3'b111;
      // memory_array[17572] <= 3'b000;
      // memory_array[17573] <= 3'b000;
      // memory_array[17574] <= 3'b111;
      // memory_array[17575] <= 3'b111;
      // memory_array[17576] <= 3'b111;
      // memory_array[17577] <= 3'b111;
      // memory_array[17578] <= 3'b111;
      // memory_array[17579] <= 3'b110;
      // memory_array[17580] <= 3'b110;
      // memory_array[17581] <= 3'b110;
      // memory_array[17582] <= 3'b110;
      // memory_array[17583] <= 3'b110;
      // memory_array[17584] <= 3'b110;
      // memory_array[17585] <= 3'b111;
      // memory_array[17586] <= 3'b111;
      // memory_array[17587] <= 3'b111;
      // memory_array[17588] <= 3'b110;
      // memory_array[17589] <= 3'b000;
      // memory_array[17590] <= 3'b000;
      // memory_array[17591] <= 3'b101;
      // memory_array[17592] <= 3'b101;
      // memory_array[17593] <= 3'b101;
      // memory_array[17594] <= 3'b101;
      // memory_array[17595] <= 3'b111;
      // memory_array[17596] <= 3'b111;
      // memory_array[17597] <= 3'b101;
      // memory_array[17598] <= 3'b101;
      // memory_array[17599] <= 3'b101;
      // memory_array[17600] <= 3'b101;
      // memory_array[17601] <= 3'b101;
      // memory_array[17602] <= 3'b101;
      // memory_array[17603] <= 3'b101;
      // memory_array[17604] <= 3'b101;
      // memory_array[17605] <= 3'b101;
      // memory_array[17606] <= 3'b101;
      // memory_array[17607] <= 3'b101;
      // memory_array[17608] <= 3'b101;
      // memory_array[17609] <= 3'b000;
      // memory_array[17610] <= 3'b000;
      // memory_array[17611] <= 3'b110;
      // memory_array[17612] <= 3'b110;
      // memory_array[17613] <= 3'b111;
      // memory_array[17614] <= 3'b111;
      // memory_array[17615] <= 3'b110;
      // memory_array[17616] <= 3'b110;
      // memory_array[17617] <= 3'b110;
      // memory_array[17618] <= 3'b111;
      // memory_array[17619] <= 3'b111;
      // memory_array[17620] <= 3'b110;
      // memory_array[17621] <= 3'b000;
      // memory_array[17622] <= 3'b110;
      // memory_array[17623] <= 3'b000;
      // memory_array[17624] <= 3'b111;
      // memory_array[17625] <= 3'b111;
      // memory_array[17626] <= 3'b111;
      // memory_array[17627] <= 3'b111;
      // memory_array[17628] <= 3'b000;
      // memory_array[17629] <= 3'b111;
      // memory_array[17630] <= 3'b110;
      // memory_array[17631] <= 3'b110;
      // memory_array[17632] <= 3'b111;
      // memory_array[17633] <= 3'b111;
      // memory_array[17634] <= 3'b111;
      // memory_array[17635] <= 3'b111;
      // memory_array[17636] <= 3'b000;
      // memory_array[17637] <= 3'b111;
      // memory_array[17638] <= 3'b111;
      // memory_array[17639] <= 3'b111;
      // memory_array[17640] <= 3'b111;
      // memory_array[17641] <= 3'b111;
      // memory_array[17642] <= 3'b000;
      // memory_array[17643] <= 3'b000;
      // memory_array[17644] <= 3'b000;
      // memory_array[17645] <= 3'b111;
      // memory_array[17646] <= 3'b111;
      // memory_array[17647] <= 3'b111;
      // memory_array[17648] <= 3'b111;
      // memory_array[17649] <= 3'b000;
      // memory_array[17650] <= 3'b000;
      // memory_array[17651] <= 3'b111;
      // memory_array[17652] <= 3'b111;
      // memory_array[17653] <= 3'b111;
      // memory_array[17654] <= 3'b111;
      // memory_array[17655] <= 3'b000;
      // memory_array[17656] <= 3'b000;
      // memory_array[17657] <= 3'b111;
      // memory_array[17658] <= 3'b111;
      // memory_array[17659] <= 3'b111;
      // memory_array[17660] <= 3'b111;
      // memory_array[17661] <= 3'b111;
      // memory_array[17662] <= 3'b000;
      // memory_array[17663] <= 3'b000;
      // memory_array[17664] <= 3'b000;
      // memory_array[17665] <= 3'b101;
      // memory_array[17666] <= 3'b000;
      // memory_array[17667] <= 3'b111;
      // memory_array[17668] <= 3'b111;
      // memory_array[17669] <= 3'b111;
      // memory_array[17670] <= 3'b111;
      // memory_array[17671] <= 3'b000;
      // memory_array[17672] <= 3'b111;
      // memory_array[17673] <= 3'b111;
      // memory_array[17674] <= 3'b111;
      // memory_array[17675] <= 3'b111;
      // memory_array[17676] <= 3'b000;
      // memory_array[17677] <= 3'b101;
      // memory_array[17678] <= 3'b000;
      // memory_array[17679] <= 3'b000;
      // memory_array[17680] <= 3'b101;
      // memory_array[17681] <= 3'b110;
      // memory_array[17682] <= 3'b000;
      // memory_array[17683] <= 3'b111;
      // memory_array[17684] <= 3'b111;
      // memory_array[17685] <= 3'b111;
      // memory_array[17686] <= 3'b111;
      // memory_array[17687] <= 3'b000;
      // memory_array[17688] <= 3'b000;
      // memory_array[17689] <= 3'b000;
      // memory_array[17690] <= 3'b000;
      // memory_array[17691] <= 3'b000;
      // memory_array[17692] <= 3'b000;
      // memory_array[17693] <= 3'b000;
      // memory_array[17694] <= 3'b000;
      // memory_array[17695] <= 3'b000;
      // memory_array[17696] <= 3'b110;
      // memory_array[17697] <= 3'b110;
      // memory_array[17698] <= 3'b110;
      // memory_array[17699] <= 3'b110;
      // memory_array[17700] <= 3'b110;
      // memory_array[17701] <= 3'b000;
      // memory_array[17702] <= 3'b111;
      // memory_array[17703] <= 3'b111;
      // memory_array[17704] <= 3'b000;
      // memory_array[17705] <= 3'b000;
      // memory_array[17706] <= 3'b000;
      // memory_array[17707] <= 3'b000;
      // memory_array[17708] <= 3'b111;
      // memory_array[17709] <= 3'b111;
      // memory_array[17710] <= 3'b111;
      // memory_array[17711] <= 3'b111;
      // memory_array[17712] <= 3'b000;
      // memory_array[17713] <= 3'b000;
      // memory_array[17714] <= 3'b000;
      // memory_array[17715] <= 3'b000;
      // memory_array[17716] <= 3'b000;
      // memory_array[17717] <= 3'b111;
      // memory_array[17718] <= 3'b111;
      // memory_array[17719] <= 3'b111;
      // memory_array[17720] <= 3'b111;
      // memory_array[17721] <= 3'b000;
      // memory_array[17722] <= 3'b111;
      // memory_array[17723] <= 3'b111;
      // memory_array[17724] <= 3'b111;
      // memory_array[17725] <= 3'b111;
      // memory_array[17726] <= 3'b000;
      // memory_array[17727] <= 3'b000;
      // memory_array[17728] <= 3'b000;
      // memory_array[17729] <= 3'b000;
      // memory_array[17730] <= 3'b000;
      // memory_array[17731] <= 3'b000;
      // memory_array[17732] <= 3'b110;
      // memory_array[17733] <= 3'b000;
      // memory_array[17734] <= 3'b000;
      // memory_array[17735] <= 3'b111;
      // memory_array[17736] <= 3'b111;
      // memory_array[17737] <= 3'b111;
      // memory_array[17738] <= 3'b111;
      // memory_array[17739] <= 3'b000;
      // memory_array[17740] <= 3'b000;
      // memory_array[17741] <= 3'b000;
      // memory_array[17742] <= 3'b000;
      // memory_array[17743] <= 3'b111;
      // memory_array[17744] <= 3'b111;
      // memory_array[17745] <= 3'b111;
      // memory_array[17746] <= 3'b111;
      // memory_array[17747] <= 3'b000;
      // memory_array[17748] <= 3'b111;
      // memory_array[17749] <= 3'b111;
      // memory_array[17750] <= 3'b111;
      // memory_array[17751] <= 3'b111;
      // memory_array[17752] <= 3'b000;
      // memory_array[17753] <= 3'b111;
      // memory_array[17754] <= 3'b000;
      // memory_array[17755] <= 3'b000;
      // memory_array[17756] <= 3'b000;
      // memory_array[17757] <= 3'b000;
      // memory_array[17758] <= 3'b000;
      // memory_array[17759] <= 3'b000;
      // memory_array[17760] <= 3'b000;
      // memory_array[17761] <= 3'b000;
      // memory_array[17762] <= 3'b111;
      // memory_array[17763] <= 3'b111;
      // memory_array[17764] <= 3'b111;
      // memory_array[17765] <= 3'b111;
      // memory_array[17766] <= 3'b110;
      // memory_array[17767] <= 3'b111;
      // memory_array[17768] <= 3'b111;
      // memory_array[17769] <= 3'b111;
      // memory_array[17770] <= 3'b111;
      // memory_array[17771] <= 3'b111;
      // memory_array[17772] <= 3'b000;
      // memory_array[17773] <= 3'b000;
      // memory_array[17774] <= 3'b111;
      // memory_array[17775] <= 3'b111;
      // memory_array[17776] <= 3'b111;
      // memory_array[17777] <= 3'b111;
      // memory_array[17778] <= 3'b111;
      // memory_array[17779] <= 3'b110;
      // memory_array[17780] <= 3'b110;
      // memory_array[17781] <= 3'b110;
      // memory_array[17782] <= 3'b110;
      // memory_array[17783] <= 3'b110;
      // memory_array[17784] <= 3'b110;
      // memory_array[17785] <= 3'b110;
      // memory_array[17786] <= 3'b110;
      // memory_array[17787] <= 3'b110;
      // memory_array[17788] <= 3'b110;
      // memory_array[17789] <= 3'b000;
      // memory_array[17790] <= 3'b000;
      // memory_array[17791] <= 3'b101;
      // memory_array[17792] <= 3'b101;
      // memory_array[17793] <= 3'b101;
      // memory_array[17794] <= 3'b101;
      // memory_array[17795] <= 3'b101;
      // memory_array[17796] <= 3'b101;
      // memory_array[17797] <= 3'b101;
      // memory_array[17798] <= 3'b101;
      // memory_array[17799] <= 3'b101;
      // memory_array[17800] <= 3'b101;
      // memory_array[17801] <= 3'b101;
      // memory_array[17802] <= 3'b101;
      // memory_array[17803] <= 3'b101;
      // memory_array[17804] <= 3'b101;
      // memory_array[17805] <= 3'b101;
      // memory_array[17806] <= 3'b101;
      // memory_array[17807] <= 3'b101;
      // memory_array[17808] <= 3'b101;
      // memory_array[17809] <= 3'b000;
      // memory_array[17810] <= 3'b000;
      // memory_array[17811] <= 3'b110;
      // memory_array[17812] <= 3'b110;
      // memory_array[17813] <= 3'b111;
      // memory_array[17814] <= 3'b111;
      // memory_array[17815] <= 3'b110;
      // memory_array[17816] <= 3'b110;
      // memory_array[17817] <= 3'b110;
      // memory_array[17818] <= 3'b111;
      // memory_array[17819] <= 3'b111;
      // memory_array[17820] <= 3'b110;
      // memory_array[17821] <= 3'b000;
      // memory_array[17822] <= 3'b110;
      // memory_array[17823] <= 3'b000;
      // memory_array[17824] <= 3'b111;
      // memory_array[17825] <= 3'b111;
      // memory_array[17826] <= 3'b111;
      // memory_array[17827] <= 3'b000;
      // memory_array[17828] <= 3'b111;
      // memory_array[17829] <= 3'b111;
      // memory_array[17830] <= 3'b110;
      // memory_array[17831] <= 3'b110;
      // memory_array[17832] <= 3'b000;
      // memory_array[17833] <= 3'b111;
      // memory_array[17834] <= 3'b111;
      // memory_array[17835] <= 3'b111;
      // memory_array[17836] <= 3'b000;
      // memory_array[17837] <= 3'b111;
      // memory_array[17838] <= 3'b111;
      // memory_array[17839] <= 3'b111;
      // memory_array[17840] <= 3'b111;
      // memory_array[17841] <= 3'b000;
      // memory_array[17842] <= 3'b000;
      // memory_array[17843] <= 3'b000;
      // memory_array[17844] <= 3'b110;
      // memory_array[17845] <= 3'b000;
      // memory_array[17846] <= 3'b111;
      // memory_array[17847] <= 3'b111;
      // memory_array[17848] <= 3'b111;
      // memory_array[17849] <= 3'b000;
      // memory_array[17850] <= 3'b000;
      // memory_array[17851] <= 3'b111;
      // memory_array[17852] <= 3'b111;
      // memory_array[17853] <= 3'b111;
      // memory_array[17854] <= 3'b111;
      // memory_array[17855] <= 3'b000;
      // memory_array[17856] <= 3'b101;
      // memory_array[17857] <= 3'b111;
      // memory_array[17858] <= 3'b111;
      // memory_array[17859] <= 3'b111;
      // memory_array[17860] <= 3'b111;
      // memory_array[17861] <= 3'b000;
      // memory_array[17862] <= 3'b101;
      // memory_array[17863] <= 3'b000;
      // memory_array[17864] <= 3'b000;
      // memory_array[17865] <= 3'b101;
      // memory_array[17866] <= 3'b101;
      // memory_array[17867] <= 3'b111;
      // memory_array[17868] <= 3'b111;
      // memory_array[17869] <= 3'b111;
      // memory_array[17870] <= 3'b111;
      // memory_array[17871] <= 3'b000;
      // memory_array[17872] <= 3'b111;
      // memory_array[17873] <= 3'b111;
      // memory_array[17874] <= 3'b111;
      // memory_array[17875] <= 3'b111;
      // memory_array[17876] <= 3'b000;
      // memory_array[17877] <= 3'b000;
      // memory_array[17878] <= 3'b000;
      // memory_array[17879] <= 3'b000;
      // memory_array[17880] <= 3'b000;
      // memory_array[17881] <= 3'b101;
      // memory_array[17882] <= 3'b000;
      // memory_array[17883] <= 3'b111;
      // memory_array[17884] <= 3'b111;
      // memory_array[17885] <= 3'b111;
      // memory_array[17886] <= 3'b000;
      // memory_array[17887] <= 3'b000;
      // memory_array[17888] <= 3'b000;
      // memory_array[17889] <= 3'b000;
      // memory_array[17890] <= 3'b000;
      // memory_array[17891] <= 3'b101;
      // memory_array[17892] <= 3'b000;
      // memory_array[17893] <= 3'b000;
      // memory_array[17894] <= 3'b000;
      // memory_array[17895] <= 3'b000;
      // memory_array[17896] <= 3'b110;
      // memory_array[17897] <= 3'b101;
      // memory_array[17898] <= 3'b000;
      // memory_array[17899] <= 3'b000;
      // memory_array[17900] <= 3'b101;
      // memory_array[17901] <= 3'b111;
      // memory_array[17902] <= 3'b111;
      // memory_array[17903] <= 3'b111;
      // memory_array[17904] <= 3'b000;
      // memory_array[17905] <= 3'b000;
      // memory_array[17906] <= 3'b101;
      // memory_array[17907] <= 3'b000;
      // memory_array[17908] <= 3'b111;
      // memory_array[17909] <= 3'b111;
      // memory_array[17910] <= 3'b111;
      // memory_array[17911] <= 3'b111;
      // memory_array[17912] <= 3'b000;
      // memory_array[17913] <= 3'b000;
      // memory_array[17914] <= 3'b000;
      // memory_array[17915] <= 3'b000;
      // memory_array[17916] <= 3'b000;
      // memory_array[17917] <= 3'b111;
      // memory_array[17918] <= 3'b111;
      // memory_array[17919] <= 3'b111;
      // memory_array[17920] <= 3'b111;
      // memory_array[17921] <= 3'b111;
      // memory_array[17922] <= 3'b111;
      // memory_array[17923] <= 3'b111;
      // memory_array[17924] <= 3'b111;
      // memory_array[17925] <= 3'b000;
      // memory_array[17926] <= 3'b000;
      // memory_array[17927] <= 3'b000;
      // memory_array[17928] <= 3'b000;
      // memory_array[17929] <= 3'b000;
      // memory_array[17930] <= 3'b000;
      // memory_array[17931] <= 3'b000;
      // memory_array[17932] <= 3'b000;
      // memory_array[17933] <= 3'b000;
      // memory_array[17934] <= 3'b000;
      // memory_array[17935] <= 3'b111;
      // memory_array[17936] <= 3'b111;
      // memory_array[17937] <= 3'b111;
      // memory_array[17938] <= 3'b111;
      // memory_array[17939] <= 3'b000;
      // memory_array[17940] <= 3'b000;
      // memory_array[17941] <= 3'b000;
      // memory_array[17942] <= 3'b000;
      // memory_array[17943] <= 3'b111;
      // memory_array[17944] <= 3'b111;
      // memory_array[17945] <= 3'b111;
      // memory_array[17946] <= 3'b111;
      // memory_array[17947] <= 3'b000;
      // memory_array[17948] <= 3'b000;
      // memory_array[17949] <= 3'b111;
      // memory_array[17950] <= 3'b111;
      // memory_array[17951] <= 3'b111;
      // memory_array[17952] <= 3'b000;
      // memory_array[17953] <= 3'b000;
      // memory_array[17954] <= 3'b000;
      // memory_array[17955] <= 3'b000;
      // memory_array[17956] <= 3'b110;
      // memory_array[17957] <= 3'b000;
      // memory_array[17958] <= 3'b000;
      // memory_array[17959] <= 3'b000;
      // memory_array[17960] <= 3'b000;
      // memory_array[17961] <= 3'b000;
      // memory_array[17962] <= 3'b111;
      // memory_array[17963] <= 3'b111;
      // memory_array[17964] <= 3'b111;
      // memory_array[17965] <= 3'b111;
      // memory_array[17966] <= 3'b110;
      // memory_array[17967] <= 3'b110;
      // memory_array[17968] <= 3'b000;
      // memory_array[17969] <= 3'b111;
      // memory_array[17970] <= 3'b111;
      // memory_array[17971] <= 3'b111;
      // memory_array[17972] <= 3'b111;
      // memory_array[17973] <= 3'b000;
      // memory_array[17974] <= 3'b000;
      // memory_array[17975] <= 3'b111;
      // memory_array[17976] <= 3'b111;
      // memory_array[17977] <= 3'b111;
      // memory_array[17978] <= 3'b111;
      // memory_array[17979] <= 3'b110;
      // memory_array[17980] <= 3'b110;
      // memory_array[17981] <= 3'b110;
      // memory_array[17982] <= 3'b110;
      // memory_array[17983] <= 3'b000;
      // memory_array[17984] <= 3'b110;
      // memory_array[17985] <= 3'b110;
      // memory_array[17986] <= 3'b110;
      // memory_array[17987] <= 3'b110;
      // memory_array[17988] <= 3'b110;
      // memory_array[17989] <= 3'b000;
      // memory_array[17990] <= 3'b000;
      // memory_array[17991] <= 3'b101;
      // memory_array[17992] <= 3'b101;
      // memory_array[17993] <= 3'b101;
      // memory_array[17994] <= 3'b101;
      // memory_array[17995] <= 3'b101;
      // memory_array[17996] <= 3'b101;
      // memory_array[17997] <= 3'b101;
      // memory_array[17998] <= 3'b101;
      // memory_array[17999] <= 3'b101;
      // memory_array[18000] <= 3'b101;
      // memory_array[18001] <= 3'b101;
      // memory_array[18002] <= 3'b101;
      // memory_array[18003] <= 3'b111;
      // memory_array[18004] <= 3'b111;
      // memory_array[18005] <= 3'b101;
      // memory_array[18006] <= 3'b101;
      // memory_array[18007] <= 3'b101;
      // memory_array[18008] <= 3'b101;
      // memory_array[18009] <= 3'b000;
      // memory_array[18010] <= 3'b000;
      // memory_array[18011] <= 3'b110;
      // memory_array[18012] <= 3'b111;
      // memory_array[18013] <= 3'b110;
      // memory_array[18014] <= 3'b110;
      // memory_array[18015] <= 3'b110;
      // memory_array[18016] <= 3'b110;
      // memory_array[18017] <= 3'b111;
      // memory_array[18018] <= 3'b110;
      // memory_array[18019] <= 3'b110;
      // memory_array[18020] <= 3'b111;
      // memory_array[18021] <= 3'b000;
      // memory_array[18022] <= 3'b110;
      // memory_array[18023] <= 3'b000;
      // memory_array[18024] <= 3'b111;
      // memory_array[18025] <= 3'b111;
      // memory_array[18026] <= 3'b111;
      // memory_array[18027] <= 3'b000;
      // memory_array[18028] <= 3'b110;
      // memory_array[18029] <= 3'b110;
      // memory_array[18030] <= 3'b111;
      // memory_array[18031] <= 3'b111;
      // memory_array[18032] <= 3'b000;
      // memory_array[18033] <= 3'b111;
      // memory_array[18034] <= 3'b111;
      // memory_array[18035] <= 3'b111;
      // memory_array[18036] <= 3'b111;
      // memory_array[18037] <= 3'b111;
      // memory_array[18038] <= 3'b111;
      // memory_array[18039] <= 3'b111;
      // memory_array[18040] <= 3'b111;
      // memory_array[18041] <= 3'b000;
      // memory_array[18042] <= 3'b000;
      // memory_array[18043] <= 3'b000;
      // memory_array[18044] <= 3'b110;
      // memory_array[18045] <= 3'b110;
      // memory_array[18046] <= 3'b111;
      // memory_array[18047] <= 3'b111;
      // memory_array[18048] <= 3'b111;
      // memory_array[18049] <= 3'b000;
      // memory_array[18050] <= 3'b000;
      // memory_array[18051] <= 3'b111;
      // memory_array[18052] <= 3'b111;
      // memory_array[18053] <= 3'b111;
      // memory_array[18054] <= 3'b111;
      // memory_array[18055] <= 3'b000;
      // memory_array[18056] <= 3'b000;
      // memory_array[18057] <= 3'b111;
      // memory_array[18058] <= 3'b111;
      // memory_array[18059] <= 3'b111;
      // memory_array[18060] <= 3'b111;
      // memory_array[18061] <= 3'b000;
      // memory_array[18062] <= 3'b101;
      // memory_array[18063] <= 3'b000;
      // memory_array[18064] <= 3'b101;
      // memory_array[18065] <= 3'b101;
      // memory_array[18066] <= 3'b000;
      // memory_array[18067] <= 3'b111;
      // memory_array[18068] <= 3'b111;
      // memory_array[18069] <= 3'b111;
      // memory_array[18070] <= 3'b111;
      // memory_array[18071] <= 3'b000;
      // memory_array[18072] <= 3'b111;
      // memory_array[18073] <= 3'b111;
      // memory_array[18074] <= 3'b111;
      // memory_array[18075] <= 3'b111;
      // memory_array[18076] <= 3'b000;
      // memory_array[18077] <= 3'b000;
      // memory_array[18078] <= 3'b000;
      // memory_array[18079] <= 3'b101;
      // memory_array[18080] <= 3'b000;
      // memory_array[18081] <= 3'b000;
      // memory_array[18082] <= 3'b111;
      // memory_array[18083] <= 3'b111;
      // memory_array[18084] <= 3'b111;
      // memory_array[18085] <= 3'b111;
      // memory_array[18086] <= 3'b000;
      // memory_array[18087] <= 3'b000;
      // memory_array[18088] <= 3'b000;
      // memory_array[18089] <= 3'b000;
      // memory_array[18090] <= 3'b000;
      // memory_array[18091] <= 3'b000;
      // memory_array[18092] <= 3'b000;
      // memory_array[18093] <= 3'b000;
      // memory_array[18094] <= 3'b111;
      // memory_array[18095] <= 3'b000;
      // memory_array[18096] <= 3'b110;
      // memory_array[18097] <= 3'b000;
      // memory_array[18098] <= 3'b101;
      // memory_array[18099] <= 3'b101;
      // memory_array[18100] <= 3'b000;
      // memory_array[18101] <= 3'b111;
      // memory_array[18102] <= 3'b111;
      // memory_array[18103] <= 3'b111;
      // memory_array[18104] <= 3'b000;
      // memory_array[18105] <= 3'b000;
      // memory_array[18106] <= 3'b000;
      // memory_array[18107] <= 3'b000;
      // memory_array[18108] <= 3'b111;
      // memory_array[18109] <= 3'b111;
      // memory_array[18110] <= 3'b111;
      // memory_array[18111] <= 3'b111;
      // memory_array[18112] <= 3'b000;
      // memory_array[18113] <= 3'b000;
      // memory_array[18114] <= 3'b000;
      // memory_array[18115] <= 3'b000;
      // memory_array[18116] <= 3'b000;
      // memory_array[18117] <= 3'b111;
      // memory_array[18118] <= 3'b111;
      // memory_array[18119] <= 3'b111;
      // memory_array[18120] <= 3'b111;
      // memory_array[18121] <= 3'b111;
      // memory_array[18122] <= 3'b111;
      // memory_array[18123] <= 3'b111;
      // memory_array[18124] <= 3'b111;
      // memory_array[18125] <= 3'b000;
      // memory_array[18126] <= 3'b000;
      // memory_array[18127] <= 3'b000;
      // memory_array[18128] <= 3'b000;
      // memory_array[18129] <= 3'b000;
      // memory_array[18130] <= 3'b000;
      // memory_array[18131] <= 3'b000;
      // memory_array[18132] <= 3'b000;
      // memory_array[18133] <= 3'b000;
      // memory_array[18134] <= 3'b000;
      // memory_array[18135] <= 3'b111;
      // memory_array[18136] <= 3'b111;
      // memory_array[18137] <= 3'b111;
      // memory_array[18138] <= 3'b111;
      // memory_array[18139] <= 3'b000;
      // memory_array[18140] <= 3'b000;
      // memory_array[18141] <= 3'b000;
      // memory_array[18142] <= 3'b000;
      // memory_array[18143] <= 3'b111;
      // memory_array[18144] <= 3'b111;
      // memory_array[18145] <= 3'b111;
      // memory_array[18146] <= 3'b111;
      // memory_array[18147] <= 3'b000;
      // memory_array[18148] <= 3'b000;
      // memory_array[18149] <= 3'b111;
      // memory_array[18150] <= 3'b111;
      // memory_array[18151] <= 3'b111;
      // memory_array[18152] <= 3'b111;
      // memory_array[18153] <= 3'b000;
      // memory_array[18154] <= 3'b110;
      // memory_array[18155] <= 3'b000;
      // memory_array[18156] <= 3'b000;
      // memory_array[18157] <= 3'b000;
      // memory_array[18158] <= 3'b000;
      // memory_array[18159] <= 3'b000;
      // memory_array[18160] <= 3'b000;
      // memory_array[18161] <= 3'b000;
      // memory_array[18162] <= 3'b111;
      // memory_array[18163] <= 3'b111;
      // memory_array[18164] <= 3'b111;
      // memory_array[18165] <= 3'b111;
      // memory_array[18166] <= 3'b110;
      // memory_array[18167] <= 3'b111;
      // memory_array[18168] <= 3'b000;
      // memory_array[18169] <= 3'b111;
      // memory_array[18170] <= 3'b111;
      // memory_array[18171] <= 3'b111;
      // memory_array[18172] <= 3'b111;
      // memory_array[18173] <= 3'b000;
      // memory_array[18174] <= 3'b000;
      // memory_array[18175] <= 3'b111;
      // memory_array[18176] <= 3'b111;
      // memory_array[18177] <= 3'b111;
      // memory_array[18178] <= 3'b111;
      // memory_array[18179] <= 3'b110;
      // memory_array[18180] <= 3'b110;
      // memory_array[18181] <= 3'b110;
      // memory_array[18182] <= 3'b110;
      // memory_array[18183] <= 3'b110;
      // memory_array[18184] <= 3'b110;
      // memory_array[18185] <= 3'b111;
      // memory_array[18186] <= 3'b111;
      // memory_array[18187] <= 3'b111;
      // memory_array[18188] <= 3'b110;
      // memory_array[18189] <= 3'b000;
      // memory_array[18190] <= 3'b000;
      // memory_array[18191] <= 3'b101;
      // memory_array[18192] <= 3'b101;
      // memory_array[18193] <= 3'b101;
      // memory_array[18194] <= 3'b101;
      // memory_array[18195] <= 3'b111;
      // memory_array[18196] <= 3'b111;
      // memory_array[18197] <= 3'b101;
      // memory_array[18198] <= 3'b101;
      // memory_array[18199] <= 3'b101;
      // memory_array[18200] <= 3'b101;
      // memory_array[18201] <= 3'b101;
      // memory_array[18202] <= 3'b110;
      // memory_array[18203] <= 3'b101;
      // memory_array[18204] <= 3'b101;
      // memory_array[18205] <= 3'b110;
      // memory_array[18206] <= 3'b101;
      // memory_array[18207] <= 3'b101;
      // memory_array[18208] <= 3'b101;
      // memory_array[18209] <= 3'b000;
      // memory_array[18210] <= 3'b000;
      // memory_array[18211] <= 3'b110;
      // memory_array[18212] <= 3'b110;
      // memory_array[18213] <= 3'b110;
      // memory_array[18214] <= 3'b110;
      // memory_array[18215] <= 3'b110;
      // memory_array[18216] <= 3'b110;
      // memory_array[18217] <= 3'b110;
      // memory_array[18218] <= 3'b110;
      // memory_array[18219] <= 3'b110;
      // memory_array[18220] <= 3'b110;
      // memory_array[18221] <= 3'b000;
      // memory_array[18222] <= 3'b110;
      // memory_array[18223] <= 3'b000;
      // memory_array[18224] <= 3'b111;
      // memory_array[18225] <= 3'b111;
      // memory_array[18226] <= 3'b111;
      // memory_array[18227] <= 3'b000;
      // memory_array[18228] <= 3'b111;
      // memory_array[18229] <= 3'b110;
      // memory_array[18230] <= 3'b110;
      // memory_array[18231] <= 3'b110;
      // memory_array[18232] <= 3'b000;
      // memory_array[18233] <= 3'b000;
      // memory_array[18234] <= 3'b111;
      // memory_array[18235] <= 3'b111;
      // memory_array[18236] <= 3'b111;
      // memory_array[18237] <= 3'b111;
      // memory_array[18238] <= 3'b111;
      // memory_array[18239] <= 3'b111;
      // memory_array[18240] <= 3'b111;
      // memory_array[18241] <= 3'b000;
      // memory_array[18242] <= 3'b000;
      // memory_array[18243] <= 3'b000;
      // memory_array[18244] <= 3'b000;
      // memory_array[18245] <= 3'b110;
      // memory_array[18246] <= 3'b111;
      // memory_array[18247] <= 3'b111;
      // memory_array[18248] <= 3'b111;
      // memory_array[18249] <= 3'b111;
      // memory_array[18250] <= 3'b000;
      // memory_array[18251] <= 3'b111;
      // memory_array[18252] <= 3'b111;
      // memory_array[18253] <= 3'b111;
      // memory_array[18254] <= 3'b111;
      // memory_array[18255] <= 3'b000;
      // memory_array[18256] <= 3'b101;
      // memory_array[18257] <= 3'b111;
      // memory_array[18258] <= 3'b111;
      // memory_array[18259] <= 3'b111;
      // memory_array[18260] <= 3'b111;
      // memory_array[18261] <= 3'b000;
      // memory_array[18262] <= 3'b101;
      // memory_array[18263] <= 3'b000;
      // memory_array[18264] <= 3'b000;
      // memory_array[18265] <= 3'b101;
      // memory_array[18266] <= 3'b000;
      // memory_array[18267] <= 3'b111;
      // memory_array[18268] <= 3'b111;
      // memory_array[18269] <= 3'b111;
      // memory_array[18270] <= 3'b111;
      // memory_array[18271] <= 3'b000;
      // memory_array[18272] <= 3'b111;
      // memory_array[18273] <= 3'b111;
      // memory_array[18274] <= 3'b111;
      // memory_array[18275] <= 3'b111;
      // memory_array[18276] <= 3'b000;
      // memory_array[18277] <= 3'b000;
      // memory_array[18278] <= 3'b000;
      // memory_array[18279] <= 3'b000;
      // memory_array[18280] <= 3'b101;
      // memory_array[18281] <= 3'b110;
      // memory_array[18282] <= 3'b111;
      // memory_array[18283] <= 3'b111;
      // memory_array[18284] <= 3'b111;
      // memory_array[18285] <= 3'b111;
      // memory_array[18286] <= 3'b000;
      // memory_array[18287] <= 3'b000;
      // memory_array[18288] <= 3'b000;
      // memory_array[18289] <= 3'b000;
      // memory_array[18290] <= 3'b000;
      // memory_array[18291] <= 3'b000;
      // memory_array[18292] <= 3'b000;
      // memory_array[18293] <= 3'b000;
      // memory_array[18294] <= 3'b111;
      // memory_array[18295] <= 3'b000;
      // memory_array[18296] <= 3'b101;
      // memory_array[18297] <= 3'b101;
      // memory_array[18298] <= 3'b000;
      // memory_array[18299] <= 3'b000;
      // memory_array[18300] <= 3'b101;
      // memory_array[18301] <= 3'b111;
      // memory_array[18302] <= 3'b111;
      // memory_array[18303] <= 3'b111;
      // memory_array[18304] <= 3'b000;
      // memory_array[18305] <= 3'b000;
      // memory_array[18306] <= 3'b101;
      // memory_array[18307] <= 3'b000;
      // memory_array[18308] <= 3'b111;
      // memory_array[18309] <= 3'b111;
      // memory_array[18310] <= 3'b111;
      // memory_array[18311] <= 3'b111;
      // memory_array[18312] <= 3'b000;
      // memory_array[18313] <= 3'b000;
      // memory_array[18314] <= 3'b000;
      // memory_array[18315] <= 3'b000;
      // memory_array[18316] <= 3'b000;
      // memory_array[18317] <= 3'b111;
      // memory_array[18318] <= 3'b111;
      // memory_array[18319] <= 3'b111;
      // memory_array[18320] <= 3'b111;
      // memory_array[18321] <= 3'b111;
      // memory_array[18322] <= 3'b111;
      // memory_array[18323] <= 3'b111;
      // memory_array[18324] <= 3'b111;
      // memory_array[18325] <= 3'b000;
      // memory_array[18326] <= 3'b000;
      // memory_array[18327] <= 3'b000;
      // memory_array[18328] <= 3'b000;
      // memory_array[18329] <= 3'b000;
      // memory_array[18330] <= 3'b000;
      // memory_array[18331] <= 3'b111;
      // memory_array[18332] <= 3'b000;
      // memory_array[18333] <= 3'b000;
      // memory_array[18334] <= 3'b000;
      // memory_array[18335] <= 3'b111;
      // memory_array[18336] <= 3'b111;
      // memory_array[18337] <= 3'b111;
      // memory_array[18338] <= 3'b111;
      // memory_array[18339] <= 3'b000;
      // memory_array[18340] <= 3'b000;
      // memory_array[18341] <= 3'b000;
      // memory_array[18342] <= 3'b000;
      // memory_array[18343] <= 3'b111;
      // memory_array[18344] <= 3'b111;
      // memory_array[18345] <= 3'b111;
      // memory_array[18346] <= 3'b111;
      // memory_array[18347] <= 3'b000;
      // memory_array[18348] <= 3'b000;
      // memory_array[18349] <= 3'b111;
      // memory_array[18350] <= 3'b111;
      // memory_array[18351] <= 3'b111;
      // memory_array[18352] <= 3'b111;
      // memory_array[18353] <= 3'b111;
      // memory_array[18354] <= 3'b110;
      // memory_array[18355] <= 3'b000;
      // memory_array[18356] <= 3'b000;
      // memory_array[18357] <= 3'b000;
      // memory_array[18358] <= 3'b000;
      // memory_array[18359] <= 3'b000;
      // memory_array[18360] <= 3'b000;
      // memory_array[18361] <= 3'b000;
      // memory_array[18362] <= 3'b111;
      // memory_array[18363] <= 3'b111;
      // memory_array[18364] <= 3'b111;
      // memory_array[18365] <= 3'b111;
      // memory_array[18366] <= 3'b110;
      // memory_array[18367] <= 3'b110;
      // memory_array[18368] <= 3'b000;
      // memory_array[18369] <= 3'b111;
      // memory_array[18370] <= 3'b111;
      // memory_array[18371] <= 3'b111;
      // memory_array[18372] <= 3'b000;
      // memory_array[18373] <= 3'b111;
      // memory_array[18374] <= 3'b000;
      // memory_array[18375] <= 3'b111;
      // memory_array[18376] <= 3'b111;
      // memory_array[18377] <= 3'b111;
      // memory_array[18378] <= 3'b111;
      // memory_array[18379] <= 3'b110;
      // memory_array[18380] <= 3'b110;
      // memory_array[18381] <= 3'b110;
      // memory_array[18382] <= 3'b110;
      // memory_array[18383] <= 3'b000;
      // memory_array[18384] <= 3'b111;
      // memory_array[18385] <= 3'b110;
      // memory_array[18386] <= 3'b110;
      // memory_array[18387] <= 3'b110;
      // memory_array[18388] <= 3'b000;
      // memory_array[18389] <= 3'b000;
      // memory_array[18390] <= 3'b000;
      // memory_array[18391] <= 3'b101;
      // memory_array[18392] <= 3'b101;
      // memory_array[18393] <= 3'b101;
      // memory_array[18394] <= 3'b000;
      // memory_array[18395] <= 3'b101;
      // memory_array[18396] <= 3'b101;
      // memory_array[18397] <= 3'b110;
      // memory_array[18398] <= 3'b101;
      // memory_array[18399] <= 3'b101;
      // memory_array[18400] <= 3'b101;
      // memory_array[18401] <= 3'b110;
      // memory_array[18402] <= 3'b110;
      // memory_array[18403] <= 3'b000;
      // memory_array[18404] <= 3'b000;
      // memory_array[18405] <= 3'b110;
      // memory_array[18406] <= 3'b110;
      // memory_array[18407] <= 3'b101;
      // memory_array[18408] <= 3'b101;
      // memory_array[18409] <= 3'b000;
      // memory_array[18410] <= 3'b000;
      // memory_array[18411] <= 3'b110;
      // memory_array[18412] <= 3'b110;
      // memory_array[18413] <= 3'b110;
      // memory_array[18414] <= 3'b110;
      // memory_array[18415] <= 3'b110;
      // memory_array[18416] <= 3'b110;
      // memory_array[18417] <= 3'b110;
      // memory_array[18418] <= 3'b111;
      // memory_array[18419] <= 3'b111;
      // memory_array[18420] <= 3'b110;
      // memory_array[18421] <= 3'b000;
      // memory_array[18422] <= 3'b110;
      // memory_array[18423] <= 3'b000;
      // memory_array[18424] <= 3'b111;
      // memory_array[18425] <= 3'b111;
      // memory_array[18426] <= 3'b111;
      // memory_array[18427] <= 3'b000;
      // memory_array[18428] <= 3'b111;
      // memory_array[18429] <= 3'b111;
      // memory_array[18430] <= 3'b110;
      // memory_array[18431] <= 3'b110;
      // memory_array[18432] <= 3'b000;
      // memory_array[18433] <= 3'b000;
      // memory_array[18434] <= 3'b111;
      // memory_array[18435] <= 3'b111;
      // memory_array[18436] <= 3'b111;
      // memory_array[18437] <= 3'b111;
      // memory_array[18438] <= 3'b111;
      // memory_array[18439] <= 3'b111;
      // memory_array[18440] <= 3'b111;
      // memory_array[18441] <= 3'b000;
      // memory_array[18442] <= 3'b110;
      // memory_array[18443] <= 3'b000;
      // memory_array[18444] <= 3'b000;
      // memory_array[18445] <= 3'b000;
      // memory_array[18446] <= 3'b111;
      // memory_array[18447] <= 3'b111;
      // memory_array[18448] <= 3'b111;
      // memory_array[18449] <= 3'b111;
      // memory_array[18450] <= 3'b000;
      // memory_array[18451] <= 3'b111;
      // memory_array[18452] <= 3'b111;
      // memory_array[18453] <= 3'b111;
      // memory_array[18454] <= 3'b111;
      // memory_array[18455] <= 3'b000;
      // memory_array[18456] <= 3'b000;
      // memory_array[18457] <= 3'b111;
      // memory_array[18458] <= 3'b111;
      // memory_array[18459] <= 3'b111;
      // memory_array[18460] <= 3'b111;
      // memory_array[18461] <= 3'b000;
      // memory_array[18462] <= 3'b101;
      // memory_array[18463] <= 3'b000;
      // memory_array[18464] <= 3'b101;
      // memory_array[18465] <= 3'b000;
      // memory_array[18466] <= 3'b000;
      // memory_array[18467] <= 3'b111;
      // memory_array[18468] <= 3'b111;
      // memory_array[18469] <= 3'b111;
      // memory_array[18470] <= 3'b111;
      // memory_array[18471] <= 3'b000;
      // memory_array[18472] <= 3'b111;
      // memory_array[18473] <= 3'b111;
      // memory_array[18474] <= 3'b111;
      // memory_array[18475] <= 3'b000;
      // memory_array[18476] <= 3'b101;
      // memory_array[18477] <= 3'b110;
      // memory_array[18478] <= 3'b000;
      // memory_array[18479] <= 3'b000;
      // memory_array[18480] <= 3'b000;
      // memory_array[18481] <= 3'b000;
      // memory_array[18482] <= 3'b111;
      // memory_array[18483] <= 3'b111;
      // memory_array[18484] <= 3'b111;
      // memory_array[18485] <= 3'b111;
      // memory_array[18486] <= 3'b000;
      // memory_array[18487] <= 3'b000;
      // memory_array[18488] <= 3'b000;
      // memory_array[18489] <= 3'b000;
      // memory_array[18490] <= 3'b000;
      // memory_array[18491] <= 3'b111;
      // memory_array[18492] <= 3'b111;
      // memory_array[18493] <= 3'b111;
      // memory_array[18494] <= 3'b000;
      // memory_array[18495] <= 3'b000;
      // memory_array[18496] <= 3'b101;
      // memory_array[18497] <= 3'b111;
      // memory_array[18498] <= 3'b111;
      // memory_array[18499] <= 3'b111;
      // memory_array[18500] <= 3'b111;
      // memory_array[18501] <= 3'b111;
      // memory_array[18502] <= 3'b111;
      // memory_array[18503] <= 3'b111;
      // memory_array[18504] <= 3'b111;
      // memory_array[18505] <= 3'b111;
      // memory_array[18506] <= 3'b000;
      // memory_array[18507] <= 3'b000;
      // memory_array[18508] <= 3'b111;
      // memory_array[18509] <= 3'b111;
      // memory_array[18510] <= 3'b111;
      // memory_array[18511] <= 3'b111;
      // memory_array[18512] <= 3'b110;
      // memory_array[18513] <= 3'b000;
      // memory_array[18514] <= 3'b000;
      // memory_array[18515] <= 3'b000;
      // memory_array[18516] <= 3'b000;
      // memory_array[18517] <= 3'b111;
      // memory_array[18518] <= 3'b111;
      // memory_array[18519] <= 3'b111;
      // memory_array[18520] <= 3'b111;
      // memory_array[18521] <= 3'b111;
      // memory_array[18522] <= 3'b111;
      // memory_array[18523] <= 3'b111;
      // memory_array[18524] <= 3'b111;
      // memory_array[18525] <= 3'b111;
      // memory_array[18526] <= 3'b111;
      // memory_array[18527] <= 3'b111;
      // memory_array[18528] <= 3'b111;
      // memory_array[18529] <= 3'b111;
      // memory_array[18530] <= 3'b111;
      // memory_array[18531] <= 3'b000;
      // memory_array[18532] <= 3'b101;
      // memory_array[18533] <= 3'b000;
      // memory_array[18534] <= 3'b000;
      // memory_array[18535] <= 3'b111;
      // memory_array[18536] <= 3'b111;
      // memory_array[18537] <= 3'b111;
      // memory_array[18538] <= 3'b111;
      // memory_array[18539] <= 3'b000;
      // memory_array[18540] <= 3'b101;
      // memory_array[18541] <= 3'b000;
      // memory_array[18542] <= 3'b000;
      // memory_array[18543] <= 3'b111;
      // memory_array[18544] <= 3'b111;
      // memory_array[18545] <= 3'b111;
      // memory_array[18546] <= 3'b111;
      // memory_array[18547] <= 3'b000;
      // memory_array[18548] <= 3'b000;
      // memory_array[18549] <= 3'b111;
      // memory_array[18550] <= 3'b111;
      // memory_array[18551] <= 3'b111;
      // memory_array[18552] <= 3'b111;
      // memory_array[18553] <= 3'b111;
      // memory_array[18554] <= 3'b000;
      // memory_array[18555] <= 3'b000;
      // memory_array[18556] <= 3'b110;
      // memory_array[18557] <= 3'b110;
      // memory_array[18558] <= 3'b110;
      // memory_array[18559] <= 3'b110;
      // memory_array[18560] <= 3'b110;
      // memory_array[18561] <= 3'b000;
      // memory_array[18562] <= 3'b111;
      // memory_array[18563] <= 3'b111;
      // memory_array[18564] <= 3'b111;
      // memory_array[18565] <= 3'b111;
      // memory_array[18566] <= 3'b110;
      // memory_array[18567] <= 3'b110;
      // memory_array[18568] <= 3'b000;
      // memory_array[18569] <= 3'b111;
      // memory_array[18570] <= 3'b111;
      // memory_array[18571] <= 3'b000;
      // memory_array[18572] <= 3'b000;
      // memory_array[18573] <= 3'b110;
      // memory_array[18574] <= 3'b000;
      // memory_array[18575] <= 3'b111;
      // memory_array[18576] <= 3'b111;
      // memory_array[18577] <= 3'b111;
      // memory_array[18578] <= 3'b111;
      // memory_array[18579] <= 3'b110;
      // memory_array[18580] <= 3'b110;
      // memory_array[18581] <= 3'b110;
      // memory_array[18582] <= 3'b110;
      // memory_array[18583] <= 3'b111;
      // memory_array[18584] <= 3'b111;
      // memory_array[18585] <= 3'b110;
      // memory_array[18586] <= 3'b110;
      // memory_array[18587] <= 3'b110;
      // memory_array[18588] <= 3'b111;
      // memory_array[18589] <= 3'b000;
      // memory_array[18590] <= 3'b000;
      // memory_array[18591] <= 3'b101;
      // memory_array[18592] <= 3'b110;
      // memory_array[18593] <= 3'b000;
      // memory_array[18594] <= 3'b000;
      // memory_array[18595] <= 3'b110;
      // memory_array[18596] <= 3'b110;
      // memory_array[18597] <= 3'b110;
      // memory_array[18598] <= 3'b000;
      // memory_array[18599] <= 3'b101;
      // memory_array[18600] <= 3'b000;
      // memory_array[18601] <= 3'b000;
      // memory_array[18602] <= 3'b000;
      // memory_array[18603] <= 3'b110;
      // memory_array[18604] <= 3'b110;
      // memory_array[18605] <= 3'b000;
      // memory_array[18606] <= 3'b000;
      // memory_array[18607] <= 3'b000;
      // memory_array[18608] <= 3'b101;
      // memory_array[18609] <= 3'b000;
      // memory_array[18610] <= 3'b000;
      // memory_array[18611] <= 3'b110;
      // memory_array[18612] <= 3'b111;
      // memory_array[18613] <= 3'b110;
      // memory_array[18614] <= 3'b110;
      // memory_array[18615] <= 3'b110;
      // memory_array[18616] <= 3'b111;
      // memory_array[18617] <= 3'b110;
      // memory_array[18618] <= 3'b110;
      // memory_array[18619] <= 3'b110;
      // memory_array[18620] <= 3'b110;
      // memory_array[18621] <= 3'b000;
      // memory_array[18622] <= 3'b111;
      // memory_array[18623] <= 3'b000;
      // memory_array[18624] <= 3'b111;
      // memory_array[18625] <= 3'b111;
      // memory_array[18626] <= 3'b111;
      // memory_array[18627] <= 3'b000;
      // memory_array[18628] <= 3'b110;
      // memory_array[18629] <= 3'b110;
      // memory_array[18630] <= 3'b110;
      // memory_array[18631] <= 3'b110;
      // memory_array[18632] <= 3'b000;
      // memory_array[18633] <= 3'b000;
      // memory_array[18634] <= 3'b111;
      // memory_array[18635] <= 3'b111;
      // memory_array[18636] <= 3'b111;
      // memory_array[18637] <= 3'b111;
      // memory_array[18638] <= 3'b111;
      // memory_array[18639] <= 3'b111;
      // memory_array[18640] <= 3'b111;
      // memory_array[18641] <= 3'b000;
      // memory_array[18642] <= 3'b000;
      // memory_array[18643] <= 3'b110;
      // memory_array[18644] <= 3'b110;
      // memory_array[18645] <= 3'b000;
      // memory_array[18646] <= 3'b111;
      // memory_array[18647] <= 3'b111;
      // memory_array[18648] <= 3'b111;
      // memory_array[18649] <= 3'b111;
      // memory_array[18650] <= 3'b000;
      // memory_array[18651] <= 3'b111;
      // memory_array[18652] <= 3'b111;
      // memory_array[18653] <= 3'b111;
      // memory_array[18654] <= 3'b111;
      // memory_array[18655] <= 3'b000;
      // memory_array[18656] <= 3'b000;
      // memory_array[18657] <= 3'b111;
      // memory_array[18658] <= 3'b111;
      // memory_array[18659] <= 3'b111;
      // memory_array[18660] <= 3'b111;
      // memory_array[18661] <= 3'b000;
      // memory_array[18662] <= 3'b000;
      // memory_array[18663] <= 3'b000;
      // memory_array[18664] <= 3'b000;
      // memory_array[18665] <= 3'b000;
      // memory_array[18666] <= 3'b000;
      // memory_array[18667] <= 3'b111;
      // memory_array[18668] <= 3'b111;
      // memory_array[18669] <= 3'b111;
      // memory_array[18670] <= 3'b111;
      // memory_array[18671] <= 3'b000;
      // memory_array[18672] <= 3'b111;
      // memory_array[18673] <= 3'b111;
      // memory_array[18674] <= 3'b111;
      // memory_array[18675] <= 3'b000;
      // memory_array[18676] <= 3'b000;
      // memory_array[18677] <= 3'b000;
      // memory_array[18678] <= 3'b101;
      // memory_array[18679] <= 3'b000;
      // memory_array[18680] <= 3'b000;
      // memory_array[18681] <= 3'b000;
      // memory_array[18682] <= 3'b111;
      // memory_array[18683] <= 3'b111;
      // memory_array[18684] <= 3'b111;
      // memory_array[18685] <= 3'b111;
      // memory_array[18686] <= 3'b111;
      // memory_array[18687] <= 3'b111;
      // memory_array[18688] <= 3'b111;
      // memory_array[18689] <= 3'b111;
      // memory_array[18690] <= 3'b111;
      // memory_array[18691] <= 3'b111;
      // memory_array[18692] <= 3'b111;
      // memory_array[18693] <= 3'b000;
      // memory_array[18694] <= 3'b000;
      // memory_array[18695] <= 3'b000;
      // memory_array[18696] <= 3'b000;
      // memory_array[18697] <= 3'b000;
      // memory_array[18698] <= 3'b111;
      // memory_array[18699] <= 3'b111;
      // memory_array[18700] <= 3'b111;
      // memory_array[18701] <= 3'b111;
      // memory_array[18702] <= 3'b111;
      // memory_array[18703] <= 3'b111;
      // memory_array[18704] <= 3'b111;
      // memory_array[18705] <= 3'b111;
      // memory_array[18706] <= 3'b000;
      // memory_array[18707] <= 3'b000;
      // memory_array[18708] <= 3'b111;
      // memory_array[18709] <= 3'b111;
      // memory_array[18710] <= 3'b111;
      // memory_array[18711] <= 3'b111;
      // memory_array[18712] <= 3'b000;
      // memory_array[18713] <= 3'b000;
      // memory_array[18714] <= 3'b000;
      // memory_array[18715] <= 3'b000;
      // memory_array[18716] <= 3'b000;
      // memory_array[18717] <= 3'b111;
      // memory_array[18718] <= 3'b111;
      // memory_array[18719] <= 3'b111;
      // memory_array[18720] <= 3'b111;
      // memory_array[18721] <= 3'b111;
      // memory_array[18722] <= 3'b111;
      // memory_array[18723] <= 3'b111;
      // memory_array[18724] <= 3'b111;
      // memory_array[18725] <= 3'b111;
      // memory_array[18726] <= 3'b111;
      // memory_array[18727] <= 3'b111;
      // memory_array[18728] <= 3'b111;
      // memory_array[18729] <= 3'b111;
      // memory_array[18730] <= 3'b111;
      // memory_array[18731] <= 3'b000;
      // memory_array[18732] <= 3'b000;
      // memory_array[18733] <= 3'b000;
      // memory_array[18734] <= 3'b000;
      // memory_array[18735] <= 3'b111;
      // memory_array[18736] <= 3'b111;
      // memory_array[18737] <= 3'b111;
      // memory_array[18738] <= 3'b111;
      // memory_array[18739] <= 3'b101;
      // memory_array[18740] <= 3'b000;
      // memory_array[18741] <= 3'b000;
      // memory_array[18742] <= 3'b000;
      // memory_array[18743] <= 3'b111;
      // memory_array[18744] <= 3'b111;
      // memory_array[18745] <= 3'b111;
      // memory_array[18746] <= 3'b111;
      // memory_array[18747] <= 3'b000;
      // memory_array[18748] <= 3'b101;
      // memory_array[18749] <= 3'b000;
      // memory_array[18750] <= 3'b111;
      // memory_array[18751] <= 3'b111;
      // memory_array[18752] <= 3'b111;
      // memory_array[18753] <= 3'b111;
      // memory_array[18754] <= 3'b111;
      // memory_array[18755] <= 3'b000;
      // memory_array[18756] <= 3'b110;
      // memory_array[18757] <= 3'b000;
      // memory_array[18758] <= 3'b110;
      // memory_array[18759] <= 3'b110;
      // memory_array[18760] <= 3'b000;
      // memory_array[18761] <= 3'b000;
      // memory_array[18762] <= 3'b111;
      // memory_array[18763] <= 3'b111;
      // memory_array[18764] <= 3'b111;
      // memory_array[18765] <= 3'b111;
      // memory_array[18766] <= 3'b110;
      // memory_array[18767] <= 3'b110;
      // memory_array[18768] <= 3'b000;
      // memory_array[18769] <= 3'b111;
      // memory_array[18770] <= 3'b111;
      // memory_array[18771] <= 3'b111;
      // memory_array[18772] <= 3'b000;
      // memory_array[18773] <= 3'b110;
      // memory_array[18774] <= 3'b000;
      // memory_array[18775] <= 3'b111;
      // memory_array[18776] <= 3'b111;
      // memory_array[18777] <= 3'b111;
      // memory_array[18778] <= 3'b111;
      // memory_array[18779] <= 3'b110;
      // memory_array[18780] <= 3'b111;
      // memory_array[18781] <= 3'b111;
      // memory_array[18782] <= 3'b111;
      // memory_array[18783] <= 3'b110;
      // memory_array[18784] <= 3'b110;
      // memory_array[18785] <= 3'b111;
      // memory_array[18786] <= 3'b111;
      // memory_array[18787] <= 3'b111;
      // memory_array[18788] <= 3'b110;
      // memory_array[18789] <= 3'b000;
      // memory_array[18790] <= 3'b000;
      // memory_array[18791] <= 3'b101;
      // memory_array[18792] <= 3'b000;
      // memory_array[18793] <= 3'b110;
      // memory_array[18794] <= 3'b110;
      // memory_array[18795] <= 3'b000;
      // memory_array[18796] <= 3'b000;
      // memory_array[18797] <= 3'b000;
      // memory_array[18798] <= 3'b110;
      // memory_array[18799] <= 3'b110;
      // memory_array[18800] <= 3'b101;
      // memory_array[18801] <= 3'b101;
      // memory_array[18802] <= 3'b101;
      // memory_array[18803] <= 3'b101;
      // memory_array[18804] <= 3'b101;
      // memory_array[18805] <= 3'b101;
      // memory_array[18806] <= 3'b101;
      // memory_array[18807] <= 3'b101;
      // memory_array[18808] <= 3'b101;
      // memory_array[18809] <= 3'b000;
      // memory_array[18810] <= 3'b000;
      // memory_array[18811] <= 3'b110;
      // memory_array[18812] <= 3'b111;
      // memory_array[18813] <= 3'b110;
      // memory_array[18814] <= 3'b110;
      // memory_array[18815] <= 3'b110;
      // memory_array[18816] <= 3'b111;
      // memory_array[18817] <= 3'b110;
      // memory_array[18818] <= 3'b110;
      // memory_array[18819] <= 3'b110;
      // memory_array[18820] <= 3'b110;
      // memory_array[18821] <= 3'b000;
      // memory_array[18822] <= 3'b111;
      // memory_array[18823] <= 3'b000;
      // memory_array[18824] <= 3'b111;
      // memory_array[18825] <= 3'b111;
      // memory_array[18826] <= 3'b111;
      // memory_array[18827] <= 3'b000;
      // memory_array[18828] <= 3'b110;
      // memory_array[18829] <= 3'b110;
      // memory_array[18830] <= 3'b110;
      // memory_array[18831] <= 3'b110;
      // memory_array[18832] <= 3'b000;
      // memory_array[18833] <= 3'b000;
      // memory_array[18834] <= 3'b111;
      // memory_array[18835] <= 3'b111;
      // memory_array[18836] <= 3'b111;
      // memory_array[18837] <= 3'b111;
      // memory_array[18838] <= 3'b111;
      // memory_array[18839] <= 3'b111;
      // memory_array[18840] <= 3'b111;
      // memory_array[18841] <= 3'b000;
      // memory_array[18842] <= 3'b000;
      // memory_array[18843] <= 3'b110;
      // memory_array[18844] <= 3'b000;
      // memory_array[18845] <= 3'b111;
      // memory_array[18846] <= 3'b111;
      // memory_array[18847] <= 3'b111;
      // memory_array[18848] <= 3'b111;
      // memory_array[18849] <= 3'b111;
      // memory_array[18850] <= 3'b000;
      // memory_array[18851] <= 3'b111;
      // memory_array[18852] <= 3'b111;
      // memory_array[18853] <= 3'b111;
      // memory_array[18854] <= 3'b111;
      // memory_array[18855] <= 3'b000;
      // memory_array[18856] <= 3'b000;
      // memory_array[18857] <= 3'b111;
      // memory_array[18858] <= 3'b111;
      // memory_array[18859] <= 3'b111;
      // memory_array[18860] <= 3'b111;
      // memory_array[18861] <= 3'b000;
      // memory_array[18862] <= 3'b000;
      // memory_array[18863] <= 3'b101;
      // memory_array[18864] <= 3'b000;
      // memory_array[18865] <= 3'b000;
      // memory_array[18866] <= 3'b000;
      // memory_array[18867] <= 3'b111;
      // memory_array[18868] <= 3'b111;
      // memory_array[18869] <= 3'b111;
      // memory_array[18870] <= 3'b111;
      // memory_array[18871] <= 3'b000;
      // memory_array[18872] <= 3'b111;
      // memory_array[18873] <= 3'b111;
      // memory_array[18874] <= 3'b111;
      // memory_array[18875] <= 3'b000;
      // memory_array[18876] <= 3'b000;
      // memory_array[18877] <= 3'b000;
      // memory_array[18878] <= 3'b101;
      // memory_array[18879] <= 3'b101;
      // memory_array[18880] <= 3'b000;
      // memory_array[18881] <= 3'b000;
      // memory_array[18882] <= 3'b111;
      // memory_array[18883] <= 3'b111;
      // memory_array[18884] <= 3'b111;
      // memory_array[18885] <= 3'b111;
      // memory_array[18886] <= 3'b111;
      // memory_array[18887] <= 3'b111;
      // memory_array[18888] <= 3'b111;
      // memory_array[18889] <= 3'b111;
      // memory_array[18890] <= 3'b111;
      // memory_array[18891] <= 3'b111;
      // memory_array[18892] <= 3'b000;
      // memory_array[18893] <= 3'b000;
      // memory_array[18894] <= 3'b111;
      // memory_array[18895] <= 3'b111;
      // memory_array[18896] <= 3'b111;
      // memory_array[18897] <= 3'b111;
      // memory_array[18898] <= 3'b111;
      // memory_array[18899] <= 3'b000;
      // memory_array[18900] <= 3'b000;
      // memory_array[18901] <= 3'b111;
      // memory_array[18902] <= 3'b111;
      // memory_array[18903] <= 3'b111;
      // memory_array[18904] <= 3'b000;
      // memory_array[18905] <= 3'b000;
      // memory_array[18906] <= 3'b000;
      // memory_array[18907] <= 3'b000;
      // memory_array[18908] <= 3'b111;
      // memory_array[18909] <= 3'b111;
      // memory_array[18910] <= 3'b111;
      // memory_array[18911] <= 3'b111;
      // memory_array[18912] <= 3'b000;
      // memory_array[18913] <= 3'b101;
      // memory_array[18914] <= 3'b101;
      // memory_array[18915] <= 3'b000;
      // memory_array[18916] <= 3'b111;
      // memory_array[18917] <= 3'b111;
      // memory_array[18918] <= 3'b111;
      // memory_array[18919] <= 3'b111;
      // memory_array[18920] <= 3'b000;
      // memory_array[18921] <= 3'b111;
      // memory_array[18922] <= 3'b111;
      // memory_array[18923] <= 3'b111;
      // memory_array[18924] <= 3'b111;
      // memory_array[18925] <= 3'b111;
      // memory_array[18926] <= 3'b111;
      // memory_array[18927] <= 3'b111;
      // memory_array[18928] <= 3'b111;
      // memory_array[18929] <= 3'b000;
      // memory_array[18930] <= 3'b000;
      // memory_array[18931] <= 3'b000;
      // memory_array[18932] <= 3'b000;
      // memory_array[18933] <= 3'b101;
      // memory_array[18934] <= 3'b000;
      // memory_array[18935] <= 3'b111;
      // memory_array[18936] <= 3'b111;
      // memory_array[18937] <= 3'b111;
      // memory_array[18938] <= 3'b111;
      // memory_array[18939] <= 3'b000;
      // memory_array[18940] <= 3'b000;
      // memory_array[18941] <= 3'b000;
      // memory_array[18942] <= 3'b111;
      // memory_array[18943] <= 3'b111;
      // memory_array[18944] <= 3'b111;
      // memory_array[18945] <= 3'b111;
      // memory_array[18946] <= 3'b111;
      // memory_array[18947] <= 3'b000;
      // memory_array[18948] <= 3'b101;
      // memory_array[18949] <= 3'b000;
      // memory_array[18950] <= 3'b000;
      // memory_array[18951] <= 3'b111;
      // memory_array[18952] <= 3'b111;
      // memory_array[18953] <= 3'b111;
      // memory_array[18954] <= 3'b111;
      // memory_array[18955] <= 3'b111;
      // memory_array[18956] <= 3'b000;
      // memory_array[18957] <= 3'b000;
      // memory_array[18958] <= 3'b110;
      // memory_array[18959] <= 3'b110;
      // memory_array[18960] <= 3'b000;
      // memory_array[18961] <= 3'b000;
      // memory_array[18962] <= 3'b111;
      // memory_array[18963] <= 3'b111;
      // memory_array[18964] <= 3'b111;
      // memory_array[18965] <= 3'b111;
      // memory_array[18966] <= 3'b000;
      // memory_array[18967] <= 3'b000;
      // memory_array[18968] <= 3'b111;
      // memory_array[18969] <= 3'b000;
      // memory_array[18970] <= 3'b111;
      // memory_array[18971] <= 3'b111;
      // memory_array[18972] <= 3'b000;
      // memory_array[18973] <= 3'b110;
      // memory_array[18974] <= 3'b000;
      // memory_array[18975] <= 3'b111;
      // memory_array[18976] <= 3'b111;
      // memory_array[18977] <= 3'b111;
      // memory_array[18978] <= 3'b111;
      // memory_array[18979] <= 3'b110;
      // memory_array[18980] <= 3'b111;
      // memory_array[18981] <= 3'b111;
      // memory_array[18982] <= 3'b111;
      // memory_array[18983] <= 3'b110;
      // memory_array[18984] <= 3'b110;
      // memory_array[18985] <= 3'b111;
      // memory_array[18986] <= 3'b111;
      // memory_array[18987] <= 3'b111;
      // memory_array[18988] <= 3'b110;
      // memory_array[18989] <= 3'b000;
      // memory_array[18990] <= 3'b000;
      // memory_array[18991] <= 3'b101;
      // memory_array[18992] <= 3'b101;
      // memory_array[18993] <= 3'b101;
      // memory_array[18994] <= 3'b101;
      // memory_array[18995] <= 3'b101;
      // memory_array[18996] <= 3'b101;
      // memory_array[18997] <= 3'b101;
      // memory_array[18998] <= 3'b101;
      // memory_array[18999] <= 3'b101;
      // memory_array[19000] <= 3'b101;
      // memory_array[19001] <= 3'b101;
      // memory_array[19002] <= 3'b101;
      // memory_array[19003] <= 3'b101;
      // memory_array[19004] <= 3'b101;
      // memory_array[19005] <= 3'b101;
      // memory_array[19006] <= 3'b101;
      // memory_array[19007] <= 3'b101;
      // memory_array[19008] <= 3'b101;
      // memory_array[19009] <= 3'b000;
      // memory_array[19010] <= 3'b000;
      // memory_array[19011] <= 3'b110;
      // memory_array[19012] <= 3'b111;
      // memory_array[19013] <= 3'b110;
      // memory_array[19014] <= 3'b110;
      // memory_array[19015] <= 3'b110;
      // memory_array[19016] <= 3'b111;
      // memory_array[19017] <= 3'b110;
      // memory_array[19018] <= 3'b110;
      // memory_array[19019] <= 3'b110;
      // memory_array[19020] <= 3'b110;
      // memory_array[19021] <= 3'b000;
      // memory_array[19022] <= 3'b111;
      // memory_array[19023] <= 3'b000;
      // memory_array[19024] <= 3'b111;
      // memory_array[19025] <= 3'b111;
      // memory_array[19026] <= 3'b111;
      // memory_array[19027] <= 3'b000;
      // memory_array[19028] <= 3'b110;
      // memory_array[19029] <= 3'b110;
      // memory_array[19030] <= 3'b110;
      // memory_array[19031] <= 3'b110;
      // memory_array[19032] <= 3'b000;
      // memory_array[19033] <= 3'b000;
      // memory_array[19034] <= 3'b111;
      // memory_array[19035] <= 3'b111;
      // memory_array[19036] <= 3'b111;
      // memory_array[19037] <= 3'b111;
      // memory_array[19038] <= 3'b111;
      // memory_array[19039] <= 3'b111;
      // memory_array[19040] <= 3'b111;
      // memory_array[19041] <= 3'b000;
      // memory_array[19042] <= 3'b000;
      // memory_array[19043] <= 3'b110;
      // memory_array[19044] <= 3'b000;
      // memory_array[19045] <= 3'b111;
      // memory_array[19046] <= 3'b111;
      // memory_array[19047] <= 3'b111;
      // memory_array[19048] <= 3'b111;
      // memory_array[19049] <= 3'b111;
      // memory_array[19050] <= 3'b000;
      // memory_array[19051] <= 3'b111;
      // memory_array[19052] <= 3'b111;
      // memory_array[19053] <= 3'b111;
      // memory_array[19054] <= 3'b111;
      // memory_array[19055] <= 3'b000;
      // memory_array[19056] <= 3'b000;
      // memory_array[19057] <= 3'b111;
      // memory_array[19058] <= 3'b111;
      // memory_array[19059] <= 3'b111;
      // memory_array[19060] <= 3'b111;
      // memory_array[19061] <= 3'b000;
      // memory_array[19062] <= 3'b000;
      // memory_array[19063] <= 3'b101;
      // memory_array[19064] <= 3'b000;
      // memory_array[19065] <= 3'b000;
      // memory_array[19066] <= 3'b000;
      // memory_array[19067] <= 3'b111;
      // memory_array[19068] <= 3'b111;
      // memory_array[19069] <= 3'b111;
      // memory_array[19070] <= 3'b111;
      // memory_array[19071] <= 3'b000;
      // memory_array[19072] <= 3'b111;
      // memory_array[19073] <= 3'b111;
      // memory_array[19074] <= 3'b111;
      // memory_array[19075] <= 3'b000;
      // memory_array[19076] <= 3'b000;
      // memory_array[19077] <= 3'b000;
      // memory_array[19078] <= 3'b101;
      // memory_array[19079] <= 3'b101;
      // memory_array[19080] <= 3'b000;
      // memory_array[19081] <= 3'b000;
      // memory_array[19082] <= 3'b111;
      // memory_array[19083] <= 3'b111;
      // memory_array[19084] <= 3'b111;
      // memory_array[19085] <= 3'b111;
      // memory_array[19086] <= 3'b111;
      // memory_array[19087] <= 3'b111;
      // memory_array[19088] <= 3'b111;
      // memory_array[19089] <= 3'b111;
      // memory_array[19090] <= 3'b111;
      // memory_array[19091] <= 3'b111;
      // memory_array[19092] <= 3'b000;
      // memory_array[19093] <= 3'b000;
      // memory_array[19094] <= 3'b111;
      // memory_array[19095] <= 3'b111;
      // memory_array[19096] <= 3'b111;
      // memory_array[19097] <= 3'b111;
      // memory_array[19098] <= 3'b111;
      // memory_array[19099] <= 3'b000;
      // memory_array[19100] <= 3'b000;
      // memory_array[19101] <= 3'b111;
      // memory_array[19102] <= 3'b111;
      // memory_array[19103] <= 3'b111;
      // memory_array[19104] <= 3'b000;
      // memory_array[19105] <= 3'b000;
      // memory_array[19106] <= 3'b000;
      // memory_array[19107] <= 3'b000;
      // memory_array[19108] <= 3'b111;
      // memory_array[19109] <= 3'b111;
      // memory_array[19110] <= 3'b111;
      // memory_array[19111] <= 3'b111;
      // memory_array[19112] <= 3'b000;
      // memory_array[19113] <= 3'b101;
      // memory_array[19114] <= 3'b101;
      // memory_array[19115] <= 3'b000;
      // memory_array[19116] <= 3'b111;
      // memory_array[19117] <= 3'b111;
      // memory_array[19118] <= 3'b111;
      // memory_array[19119] <= 3'b111;
      // memory_array[19120] <= 3'b000;
      // memory_array[19121] <= 3'b111;
      // memory_array[19122] <= 3'b111;
      // memory_array[19123] <= 3'b111;
      // memory_array[19124] <= 3'b111;
      // memory_array[19125] <= 3'b111;
      // memory_array[19126] <= 3'b111;
      // memory_array[19127] <= 3'b111;
      // memory_array[19128] <= 3'b111;
      // memory_array[19129] <= 3'b000;
      // memory_array[19130] <= 3'b000;
      // memory_array[19131] <= 3'b000;
      // memory_array[19132] <= 3'b000;
      // memory_array[19133] <= 3'b101;
      // memory_array[19134] <= 3'b000;
      // memory_array[19135] <= 3'b111;
      // memory_array[19136] <= 3'b111;
      // memory_array[19137] <= 3'b111;
      // memory_array[19138] <= 3'b111;
      // memory_array[19139] <= 3'b000;
      // memory_array[19140] <= 3'b000;
      // memory_array[19141] <= 3'b000;
      // memory_array[19142] <= 3'b111;
      // memory_array[19143] <= 3'b111;
      // memory_array[19144] <= 3'b111;
      // memory_array[19145] <= 3'b111;
      // memory_array[19146] <= 3'b111;
      // memory_array[19147] <= 3'b000;
      // memory_array[19148] <= 3'b101;
      // memory_array[19149] <= 3'b000;
      // memory_array[19150] <= 3'b000;
      // memory_array[19151] <= 3'b111;
      // memory_array[19152] <= 3'b111;
      // memory_array[19153] <= 3'b111;
      // memory_array[19154] <= 3'b111;
      // memory_array[19155] <= 3'b111;
      // memory_array[19156] <= 3'b000;
      // memory_array[19157] <= 3'b000;
      // memory_array[19158] <= 3'b110;
      // memory_array[19159] <= 3'b110;
      // memory_array[19160] <= 3'b000;
      // memory_array[19161] <= 3'b000;
      // memory_array[19162] <= 3'b111;
      // memory_array[19163] <= 3'b111;
      // memory_array[19164] <= 3'b111;
      // memory_array[19165] <= 3'b111;
      // memory_array[19166] <= 3'b000;
      // memory_array[19167] <= 3'b000;
      // memory_array[19168] <= 3'b111;
      // memory_array[19169] <= 3'b000;
      // memory_array[19170] <= 3'b111;
      // memory_array[19171] <= 3'b111;
      // memory_array[19172] <= 3'b000;
      // memory_array[19173] <= 3'b110;
      // memory_array[19174] <= 3'b000;
      // memory_array[19175] <= 3'b111;
      // memory_array[19176] <= 3'b111;
      // memory_array[19177] <= 3'b111;
      // memory_array[19178] <= 3'b111;
      // memory_array[19179] <= 3'b110;
      // memory_array[19180] <= 3'b111;
      // memory_array[19181] <= 3'b111;
      // memory_array[19182] <= 3'b111;
      // memory_array[19183] <= 3'b110;
      // memory_array[19184] <= 3'b110;
      // memory_array[19185] <= 3'b111;
      // memory_array[19186] <= 3'b111;
      // memory_array[19187] <= 3'b111;
      // memory_array[19188] <= 3'b110;
      // memory_array[19189] <= 3'b000;
      // memory_array[19190] <= 3'b000;
      // memory_array[19191] <= 3'b101;
      // memory_array[19192] <= 3'b101;
      // memory_array[19193] <= 3'b101;
      // memory_array[19194] <= 3'b101;
      // memory_array[19195] <= 3'b101;
      // memory_array[19196] <= 3'b101;
      // memory_array[19197] <= 3'b101;
      // memory_array[19198] <= 3'b101;
      // memory_array[19199] <= 3'b101;
      // memory_array[19200] <= 3'b000;
      // memory_array[19201] <= 3'b000;
      // memory_array[19202] <= 3'b000;
      // memory_array[19203] <= 3'b110;
      // memory_array[19204] <= 3'b110;
      // memory_array[19205] <= 3'b000;
      // memory_array[19206] <= 3'b000;
      // memory_array[19207] <= 3'b000;
      // memory_array[19208] <= 3'b101;
      // memory_array[19209] <= 3'b000;
      // memory_array[19210] <= 3'b000;
      // memory_array[19211] <= 3'b110;
      // memory_array[19212] <= 3'b111;
      // memory_array[19213] <= 3'b110;
      // memory_array[19214] <= 3'b110;
      // memory_array[19215] <= 3'b110;
      // memory_array[19216] <= 3'b111;
      // memory_array[19217] <= 3'b110;
      // memory_array[19218] <= 3'b110;
      // memory_array[19219] <= 3'b110;
      // memory_array[19220] <= 3'b110;
      // memory_array[19221] <= 3'b000;
      // memory_array[19222] <= 3'b111;
      // memory_array[19223] <= 3'b000;
      // memory_array[19224] <= 3'b111;
      // memory_array[19225] <= 3'b111;
      // memory_array[19226] <= 3'b111;
      // memory_array[19227] <= 3'b000;
      // memory_array[19228] <= 3'b110;
      // memory_array[19229] <= 3'b110;
      // memory_array[19230] <= 3'b110;
      // memory_array[19231] <= 3'b110;
      // memory_array[19232] <= 3'b000;
      // memory_array[19233] <= 3'b000;
      // memory_array[19234] <= 3'b111;
      // memory_array[19235] <= 3'b111;
      // memory_array[19236] <= 3'b111;
      // memory_array[19237] <= 3'b111;
      // memory_array[19238] <= 3'b111;
      // memory_array[19239] <= 3'b111;
      // memory_array[19240] <= 3'b111;
      // memory_array[19241] <= 3'b000;
      // memory_array[19242] <= 3'b000;
      // memory_array[19243] <= 3'b110;
      // memory_array[19244] <= 3'b110;
      // memory_array[19245] <= 3'b000;
      // memory_array[19246] <= 3'b111;
      // memory_array[19247] <= 3'b111;
      // memory_array[19248] <= 3'b111;
      // memory_array[19249] <= 3'b000;
      // memory_array[19250] <= 3'b000;
      // memory_array[19251] <= 3'b111;
      // memory_array[19252] <= 3'b111;
      // memory_array[19253] <= 3'b111;
      // memory_array[19254] <= 3'b111;
      // memory_array[19255] <= 3'b000;
      // memory_array[19256] <= 3'b000;
      // memory_array[19257] <= 3'b111;
      // memory_array[19258] <= 3'b111;
      // memory_array[19259] <= 3'b111;
      // memory_array[19260] <= 3'b111;
      // memory_array[19261] <= 3'b000;
      // memory_array[19262] <= 3'b000;
      // memory_array[19263] <= 3'b000;
      // memory_array[19264] <= 3'b101;
      // memory_array[19265] <= 3'b000;
      // memory_array[19266] <= 3'b000;
      // memory_array[19267] <= 3'b111;
      // memory_array[19268] <= 3'b111;
      // memory_array[19269] <= 3'b111;
      // memory_array[19270] <= 3'b111;
      // memory_array[19271] <= 3'b000;
      // memory_array[19272] <= 3'b111;
      // memory_array[19273] <= 3'b111;
      // memory_array[19274] <= 3'b111;
      // memory_array[19275] <= 3'b000;
      // memory_array[19276] <= 3'b000;
      // memory_array[19277] <= 3'b000;
      // memory_array[19278] <= 3'b110;
      // memory_array[19279] <= 3'b101;
      // memory_array[19280] <= 3'b000;
      // memory_array[19281] <= 3'b000;
      // memory_array[19282] <= 3'b111;
      // memory_array[19283] <= 3'b111;
      // memory_array[19284] <= 3'b111;
      // memory_array[19285] <= 3'b111;
      // memory_array[19286] <= 3'b000;
      // memory_array[19287] <= 3'b000;
      // memory_array[19288] <= 3'b000;
      // memory_array[19289] <= 3'b000;
      // memory_array[19290] <= 3'b111;
      // memory_array[19291] <= 3'b000;
      // memory_array[19292] <= 3'b000;
      // memory_array[19293] <= 3'b000;
      // memory_array[19294] <= 3'b111;
      // memory_array[19295] <= 3'b111;
      // memory_array[19296] <= 3'b000;
      // memory_array[19297] <= 3'b000;
      // memory_array[19298] <= 3'b111;
      // memory_array[19299] <= 3'b111;
      // memory_array[19300] <= 3'b111;
      // memory_array[19301] <= 3'b111;
      // memory_array[19302] <= 3'b111;
      // memory_array[19303] <= 3'b111;
      // memory_array[19304] <= 3'b101;
      // memory_array[19305] <= 3'b000;
      // memory_array[19306] <= 3'b000;
      // memory_array[19307] <= 3'b000;
      // memory_array[19308] <= 3'b111;
      // memory_array[19309] <= 3'b111;
      // memory_array[19310] <= 3'b111;
      // memory_array[19311] <= 3'b111;
      // memory_array[19312] <= 3'b000;
      // memory_array[19313] <= 3'b101;
      // memory_array[19314] <= 3'b000;
      // memory_array[19315] <= 3'b000;
      // memory_array[19316] <= 3'b111;
      // memory_array[19317] <= 3'b111;
      // memory_array[19318] <= 3'b111;
      // memory_array[19319] <= 3'b000;
      // memory_array[19320] <= 3'b110;
      // memory_array[19321] <= 3'b111;
      // memory_array[19322] <= 3'b111;
      // memory_array[19323] <= 3'b111;
      // memory_array[19324] <= 3'b111;
      // memory_array[19325] <= 3'b000;
      // memory_array[19326] <= 3'b000;
      // memory_array[19327] <= 3'b000;
      // memory_array[19328] <= 3'b111;
      // memory_array[19329] <= 3'b000;
      // memory_array[19330] <= 3'b000;
      // memory_array[19331] <= 3'b000;
      // memory_array[19332] <= 3'b000;
      // memory_array[19333] <= 3'b000;
      // memory_array[19334] <= 3'b000;
      // memory_array[19335] <= 3'b111;
      // memory_array[19336] <= 3'b111;
      // memory_array[19337] <= 3'b111;
      // memory_array[19338] <= 3'b111;
      // memory_array[19339] <= 3'b101;
      // memory_array[19340] <= 3'b000;
      // memory_array[19341] <= 3'b111;
      // memory_array[19342] <= 3'b111;
      // memory_array[19343] <= 3'b111;
      // memory_array[19344] <= 3'b111;
      // memory_array[19345] <= 3'b111;
      // memory_array[19346] <= 3'b000;
      // memory_array[19347] <= 3'b000;
      // memory_array[19348] <= 3'b101;
      // memory_array[19349] <= 3'b000;
      // memory_array[19350] <= 3'b000;
      // memory_array[19351] <= 3'b111;
      // memory_array[19352] <= 3'b111;
      // memory_array[19353] <= 3'b111;
      // memory_array[19354] <= 3'b111;
      // memory_array[19355] <= 3'b111;
      // memory_array[19356] <= 3'b111;
      // memory_array[19357] <= 3'b000;
      // memory_array[19358] <= 3'b110;
      // memory_array[19359] <= 3'b110;
      // memory_array[19360] <= 3'b000;
      // memory_array[19361] <= 3'b000;
      // memory_array[19362] <= 3'b111;
      // memory_array[19363] <= 3'b111;
      // memory_array[19364] <= 3'b111;
      // memory_array[19365] <= 3'b111;
      // memory_array[19366] <= 3'b000;
      // memory_array[19367] <= 3'b000;
      // memory_array[19368] <= 3'b111;
      // memory_array[19369] <= 3'b110;
      // memory_array[19370] <= 3'b111;
      // memory_array[19371] <= 3'b111;
      // memory_array[19372] <= 3'b000;
      // memory_array[19373] <= 3'b000;
      // memory_array[19374] <= 3'b111;
      // memory_array[19375] <= 3'b111;
      // memory_array[19376] <= 3'b111;
      // memory_array[19377] <= 3'b111;
      // memory_array[19378] <= 3'b111;
      // memory_array[19379] <= 3'b110;
      // memory_array[19380] <= 3'b111;
      // memory_array[19381] <= 3'b111;
      // memory_array[19382] <= 3'b111;
      // memory_array[19383] <= 3'b110;
      // memory_array[19384] <= 3'b110;
      // memory_array[19385] <= 3'b111;
      // memory_array[19386] <= 3'b111;
      // memory_array[19387] <= 3'b111;
      // memory_array[19388] <= 3'b110;
      // memory_array[19389] <= 3'b000;
      // memory_array[19390] <= 3'b000;
      // memory_array[19391] <= 3'b101;
      // memory_array[19392] <= 3'b000;
      // memory_array[19393] <= 3'b110;
      // memory_array[19394] <= 3'b110;
      // memory_array[19395] <= 3'b000;
      // memory_array[19396] <= 3'b000;
      // memory_array[19397] <= 3'b000;
      // memory_array[19398] <= 3'b110;
      // memory_array[19399] <= 3'b110;
      // memory_array[19400] <= 3'b101;
      // memory_array[19401] <= 3'b000;
      // memory_array[19402] <= 3'b000;
      // memory_array[19403] <= 3'b110;
      // memory_array[19404] <= 3'b110;
      // memory_array[19405] <= 3'b000;
      // memory_array[19406] <= 3'b000;
      // memory_array[19407] <= 3'b101;
      // memory_array[19408] <= 3'b101;
      // memory_array[19409] <= 3'b000;
      // memory_array[19410] <= 3'b000;
      // memory_array[19411] <= 3'b000;
      // memory_array[19412] <= 3'b000;
      // memory_array[19413] <= 3'b000;
      // memory_array[19414] <= 3'b000;
      // memory_array[19415] <= 3'b000;
      // memory_array[19416] <= 3'b000;
      // memory_array[19417] <= 3'b000;
      // memory_array[19418] <= 3'b000;
      // memory_array[19419] <= 3'b000;
      // memory_array[19420] <= 3'b000;
      // memory_array[19421] <= 3'b000;
      // memory_array[19422] <= 3'b000;
      // memory_array[19423] <= 3'b000;
      // memory_array[19424] <= 3'b111;
      // memory_array[19425] <= 3'b111;
      // memory_array[19426] <= 3'b111;
      // memory_array[19427] <= 3'b000;
      // memory_array[19428] <= 3'b000;
      // memory_array[19429] <= 3'b000;
      // memory_array[19430] <= 3'b000;
      // memory_array[19431] <= 3'b000;
      // memory_array[19432] <= 3'b000;
      // memory_array[19433] <= 3'b000;
      // memory_array[19434] <= 3'b111;
      // memory_array[19435] <= 3'b111;
      // memory_array[19436] <= 3'b111;
      // memory_array[19437] <= 3'b111;
      // memory_array[19438] <= 3'b111;
      // memory_array[19439] <= 3'b111;
      // memory_array[19440] <= 3'b111;
      // memory_array[19441] <= 3'b000;
      // memory_array[19442] <= 3'b000;
      // memory_array[19443] <= 3'b000;
      // memory_array[19444] <= 3'b111;
      // memory_array[19445] <= 3'b000;
      // memory_array[19446] <= 3'b111;
      // memory_array[19447] <= 3'b111;
      // memory_array[19448] <= 3'b111;
      // memory_array[19449] <= 3'b000;
      // memory_array[19450] <= 3'b000;
      // memory_array[19451] <= 3'b111;
      // memory_array[19452] <= 3'b111;
      // memory_array[19453] <= 3'b111;
      // memory_array[19454] <= 3'b111;
      // memory_array[19455] <= 3'b000;
      // memory_array[19456] <= 3'b000;
      // memory_array[19457] <= 3'b111;
      // memory_array[19458] <= 3'b111;
      // memory_array[19459] <= 3'b111;
      // memory_array[19460] <= 3'b111;
      // memory_array[19461] <= 3'b000;
      // memory_array[19462] <= 3'b000;
      // memory_array[19463] <= 3'b101;
      // memory_array[19464] <= 3'b000;
      // memory_array[19465] <= 3'b000;
      // memory_array[19466] <= 3'b000;
      // memory_array[19467] <= 3'b111;
      // memory_array[19468] <= 3'b111;
      // memory_array[19469] <= 3'b111;
      // memory_array[19470] <= 3'b111;
      // memory_array[19471] <= 3'b000;
      // memory_array[19472] <= 3'b111;
      // memory_array[19473] <= 3'b111;
      // memory_array[19474] <= 3'b111;
      // memory_array[19475] <= 3'b111;
      // memory_array[19476] <= 3'b000;
      // memory_array[19477] <= 3'b000;
      // memory_array[19478] <= 3'b000;
      // memory_array[19479] <= 3'b101;
      // memory_array[19480] <= 3'b000;
      // memory_array[19481] <= 3'b000;
      // memory_array[19482] <= 3'b111;
      // memory_array[19483] <= 3'b111;
      // memory_array[19484] <= 3'b111;
      // memory_array[19485] <= 3'b111;
      // memory_array[19486] <= 3'b000;
      // memory_array[19487] <= 3'b000;
      // memory_array[19488] <= 3'b000;
      // memory_array[19489] <= 3'b000;
      // memory_array[19490] <= 3'b000;
      // memory_array[19491] <= 3'b000;
      // memory_array[19492] <= 3'b000;
      // memory_array[19493] <= 3'b000;
      // memory_array[19494] <= 3'b111;
      // memory_array[19495] <= 3'b111;
      // memory_array[19496] <= 3'b111;
      // memory_array[19497] <= 3'b000;
      // memory_array[19498] <= 3'b111;
      // memory_array[19499] <= 3'b111;
      // memory_array[19500] <= 3'b111;
      // memory_array[19501] <= 3'b111;
      // memory_array[19502] <= 3'b111;
      // memory_array[19503] <= 3'b111;
      // memory_array[19504] <= 3'b101;
      // memory_array[19505] <= 3'b000;
      // memory_array[19506] <= 3'b000;
      // memory_array[19507] <= 3'b000;
      // memory_array[19508] <= 3'b111;
      // memory_array[19509] <= 3'b111;
      // memory_array[19510] <= 3'b111;
      // memory_array[19511] <= 3'b111;
      // memory_array[19512] <= 3'b111;
      // memory_array[19513] <= 3'b111;
      // memory_array[19514] <= 3'b111;
      // memory_array[19515] <= 3'b111;
      // memory_array[19516] <= 3'b111;
      // memory_array[19517] <= 3'b000;
      // memory_array[19518] <= 3'b101;
      // memory_array[19519] <= 3'b101;
      // memory_array[19520] <= 3'b000;
      // memory_array[19521] <= 3'b111;
      // memory_array[19522] <= 3'b111;
      // memory_array[19523] <= 3'b111;
      // memory_array[19524] <= 3'b111;
      // memory_array[19525] <= 3'b000;
      // memory_array[19526] <= 3'b000;
      // memory_array[19527] <= 3'b000;
      // memory_array[19528] <= 3'b000;
      // memory_array[19529] <= 3'b101;
      // memory_array[19530] <= 3'b000;
      // memory_array[19531] <= 3'b000;
      // memory_array[19532] <= 3'b000;
      // memory_array[19533] <= 3'b101;
      // memory_array[19534] <= 3'b000;
      // memory_array[19535] <= 3'b111;
      // memory_array[19536] <= 3'b111;
      // memory_array[19537] <= 3'b111;
      // memory_array[19538] <= 3'b111;
      // memory_array[19539] <= 3'b111;
      // memory_array[19540] <= 3'b111;
      // memory_array[19541] <= 3'b111;
      // memory_array[19542] <= 3'b111;
      // memory_array[19543] <= 3'b111;
      // memory_array[19544] <= 3'b000;
      // memory_array[19545] <= 3'b000;
      // memory_array[19546] <= 3'b000;
      // memory_array[19547] <= 3'b000;
      // memory_array[19548] <= 3'b000;
      // memory_array[19549] <= 3'b000;
      // memory_array[19550] <= 3'b000;
      // memory_array[19551] <= 3'b111;
      // memory_array[19552] <= 3'b111;
      // memory_array[19553] <= 3'b111;
      // memory_array[19554] <= 3'b111;
      // memory_array[19555] <= 3'b111;
      // memory_array[19556] <= 3'b111;
      // memory_array[19557] <= 3'b000;
      // memory_array[19558] <= 3'b000;
      // memory_array[19559] <= 3'b000;
      // memory_array[19560] <= 3'b000;
      // memory_array[19561] <= 3'b000;
      // memory_array[19562] <= 3'b111;
      // memory_array[19563] <= 3'b111;
      // memory_array[19564] <= 3'b111;
      // memory_array[19565] <= 3'b111;
      // memory_array[19566] <= 3'b000;
      // memory_array[19567] <= 3'b000;
      // memory_array[19568] <= 3'b000;
      // memory_array[19569] <= 3'b000;
      // memory_array[19570] <= 3'b000;
      // memory_array[19571] <= 3'b000;
      // memory_array[19572] <= 3'b111;
      // memory_array[19573] <= 3'b111;
      // memory_array[19574] <= 3'b111;
      // memory_array[19575] <= 3'b111;
      // memory_array[19576] <= 3'b111;
      // memory_array[19577] <= 3'b111;
      // memory_array[19578] <= 3'b111;
      // memory_array[19579] <= 3'b000;
      // memory_array[19580] <= 3'b000;
      // memory_array[19581] <= 3'b000;
      // memory_array[19582] <= 3'b000;
      // memory_array[19583] <= 3'b000;
      // memory_array[19584] <= 3'b000;
      // memory_array[19585] <= 3'b000;
      // memory_array[19586] <= 3'b000;
      // memory_array[19587] <= 3'b000;
      // memory_array[19588] <= 3'b000;
      // memory_array[19589] <= 3'b000;
      // memory_array[19590] <= 3'b000;
      // memory_array[19591] <= 3'b101;
      // memory_array[19592] <= 3'b101;
      // memory_array[19593] <= 3'b110;
      // memory_array[19594] <= 3'b110;
      // memory_array[19595] <= 3'b000;
      // memory_array[19596] <= 3'b000;
      // memory_array[19597] <= 3'b000;
      // memory_array[19598] <= 3'b110;
      // memory_array[19599] <= 3'b101;
      // memory_array[19600] <= 3'b101;
      // memory_array[19601] <= 3'b101;
      // memory_array[19602] <= 3'b110;
      // memory_array[19603] <= 3'b101;
      // memory_array[19604] <= 3'b101;
      // memory_array[19605] <= 3'b110;
      // memory_array[19606] <= 3'b101;
      // memory_array[19607] <= 3'b101;
      // memory_array[19608] <= 3'b101;
      // memory_array[19609] <= 3'b000;
      // memory_array[19610] <= 3'b000;
      // memory_array[19611] <= 3'b110;
      // memory_array[19612] <= 3'b110;
      // memory_array[19613] <= 3'b110;
      // memory_array[19614] <= 3'b110;
      // memory_array[19615] <= 3'b110;
      // memory_array[19616] <= 3'b110;
      // memory_array[19617] <= 3'b110;
      // memory_array[19618] <= 3'b110;
      // memory_array[19619] <= 3'b110;
      // memory_array[19620] <= 3'b110;
      // memory_array[19621] <= 3'b000;
      // memory_array[19622] <= 3'b110;
      // memory_array[19623] <= 3'b000;
      // memory_array[19624] <= 3'b111;
      // memory_array[19625] <= 3'b111;
      // memory_array[19626] <= 3'b111;
      // memory_array[19627] <= 3'b000;
      // memory_array[19628] <= 3'b110;
      // memory_array[19629] <= 3'b110;
      // memory_array[19630] <= 3'b110;
      // memory_array[19631] <= 3'b110;
      // memory_array[19632] <= 3'b000;
      // memory_array[19633] <= 3'b111;
      // memory_array[19634] <= 3'b111;
      // memory_array[19635] <= 3'b111;
      // memory_array[19636] <= 3'b000;
      // memory_array[19637] <= 3'b111;
      // memory_array[19638] <= 3'b111;
      // memory_array[19639] <= 3'b111;
      // memory_array[19640] <= 3'b111;
      // memory_array[19641] <= 3'b000;
      // memory_array[19642] <= 3'b110;
      // memory_array[19643] <= 3'b000;
      // memory_array[19644] <= 3'b000;
      // memory_array[19645] <= 3'b111;
      // memory_array[19646] <= 3'b111;
      // memory_array[19647] <= 3'b111;
      // memory_array[19648] <= 3'b111;
      // memory_array[19649] <= 3'b101;
      // memory_array[19650] <= 3'b000;
      // memory_array[19651] <= 3'b111;
      // memory_array[19652] <= 3'b111;
      // memory_array[19653] <= 3'b111;
      // memory_array[19654] <= 3'b111;
      // memory_array[19655] <= 3'b000;
      // memory_array[19656] <= 3'b000;
      // memory_array[19657] <= 3'b111;
      // memory_array[19658] <= 3'b111;
      // memory_array[19659] <= 3'b111;
      // memory_array[19660] <= 3'b111;
      // memory_array[19661] <= 3'b000;
      // memory_array[19662] <= 3'b101;
      // memory_array[19663] <= 3'b000;
      // memory_array[19664] <= 3'b000;
      // memory_array[19665] <= 3'b000;
      // memory_array[19666] <= 3'b000;
      // memory_array[19667] <= 3'b111;
      // memory_array[19668] <= 3'b111;
      // memory_array[19669] <= 3'b111;
      // memory_array[19670] <= 3'b111;
      // memory_array[19671] <= 3'b000;
      // memory_array[19672] <= 3'b111;
      // memory_array[19673] <= 3'b111;
      // memory_array[19674] <= 3'b111;
      // memory_array[19675] <= 3'b111;
      // memory_array[19676] <= 3'b101;
      // memory_array[19677] <= 3'b000;
      // memory_array[19678] <= 3'b000;
      // memory_array[19679] <= 3'b000;
      // memory_array[19680] <= 3'b101;
      // memory_array[19681] <= 3'b000;
      // memory_array[19682] <= 3'b111;
      // memory_array[19683] <= 3'b111;
      // memory_array[19684] <= 3'b111;
      // memory_array[19685] <= 3'b111;
      // memory_array[19686] <= 3'b000;
      // memory_array[19687] <= 3'b000;
      // memory_array[19688] <= 3'b000;
      // memory_array[19689] <= 3'b000;
      // memory_array[19690] <= 3'b101;
      // memory_array[19691] <= 3'b101;
      // memory_array[19692] <= 3'b101;
      // memory_array[19693] <= 3'b000;
      // memory_array[19694] <= 3'b111;
      // memory_array[19695] <= 3'b111;
      // memory_array[19696] <= 3'b111;
      // memory_array[19697] <= 3'b111;
      // memory_array[19698] <= 3'b111;
      // memory_array[19699] <= 3'b111;
      // memory_array[19700] <= 3'b000;
      // memory_array[19701] <= 3'b111;
      // memory_array[19702] <= 3'b111;
      // memory_array[19703] <= 3'b111;
      // memory_array[19704] <= 3'b000;
      // memory_array[19705] <= 3'b000;
      // memory_array[19706] <= 3'b101;
      // memory_array[19707] <= 3'b000;
      // memory_array[19708] <= 3'b111;
      // memory_array[19709] <= 3'b111;
      // memory_array[19710] <= 3'b111;
      // memory_array[19711] <= 3'b111;
      // memory_array[19712] <= 3'b111;
      // memory_array[19713] <= 3'b111;
      // memory_array[19714] <= 3'b111;
      // memory_array[19715] <= 3'b111;
      // memory_array[19716] <= 3'b111;
      // memory_array[19717] <= 3'b000;
      // memory_array[19718] <= 3'b000;
      // memory_array[19719] <= 3'b000;
      // memory_array[19720] <= 3'b101;
      // memory_array[19721] <= 3'b111;
      // memory_array[19722] <= 3'b111;
      // memory_array[19723] <= 3'b111;
      // memory_array[19724] <= 3'b111;
      // memory_array[19725] <= 3'b000;
      // memory_array[19726] <= 3'b101;
      // memory_array[19727] <= 3'b000;
      // memory_array[19728] <= 3'b000;
      // memory_array[19729] <= 3'b000;
      // memory_array[19730] <= 3'b000;
      // memory_array[19731] <= 3'b101;
      // memory_array[19732] <= 3'b101;
      // memory_array[19733] <= 3'b000;
      // memory_array[19734] <= 3'b000;
      // memory_array[19735] <= 3'b111;
      // memory_array[19736] <= 3'b111;
      // memory_array[19737] <= 3'b111;
      // memory_array[19738] <= 3'b111;
      // memory_array[19739] <= 3'b111;
      // memory_array[19740] <= 3'b111;
      // memory_array[19741] <= 3'b111;
      // memory_array[19742] <= 3'b111;
      // memory_array[19743] <= 3'b000;
      // memory_array[19744] <= 3'b000;
      // memory_array[19745] <= 3'b101;
      // memory_array[19746] <= 3'b000;
      // memory_array[19747] <= 3'b000;
      // memory_array[19748] <= 3'b000;
      // memory_array[19749] <= 3'b000;
      // memory_array[19750] <= 3'b111;
      // memory_array[19751] <= 3'b111;
      // memory_array[19752] <= 3'b111;
      // memory_array[19753] <= 3'b111;
      // memory_array[19754] <= 3'b111;
      // memory_array[19755] <= 3'b111;
      // memory_array[19756] <= 3'b111;
      // memory_array[19757] <= 3'b111;
      // memory_array[19758] <= 3'b000;
      // memory_array[19759] <= 3'b110;
      // memory_array[19760] <= 3'b110;
      // memory_array[19761] <= 3'b000;
      // memory_array[19762] <= 3'b111;
      // memory_array[19763] <= 3'b111;
      // memory_array[19764] <= 3'b111;
      // memory_array[19765] <= 3'b111;
      // memory_array[19766] <= 3'b110;
      // memory_array[19767] <= 3'b110;
      // memory_array[19768] <= 3'b111;
      // memory_array[19769] <= 3'b111;
      // memory_array[19770] <= 3'b110;
      // memory_array[19771] <= 3'b000;
      // memory_array[19772] <= 3'b111;
      // memory_array[19773] <= 3'b111;
      // memory_array[19774] <= 3'b111;
      // memory_array[19775] <= 3'b111;
      // memory_array[19776] <= 3'b111;
      // memory_array[19777] <= 3'b111;
      // memory_array[19778] <= 3'b111;
      // memory_array[19779] <= 3'b111;
      // memory_array[19780] <= 3'b110;
      // memory_array[19781] <= 3'b110;
      // memory_array[19782] <= 3'b110;
      // memory_array[19783] <= 3'b110;
      // memory_array[19784] <= 3'b000;
      // memory_array[19785] <= 3'b110;
      // memory_array[19786] <= 3'b110;
      // memory_array[19787] <= 3'b110;
      // memory_array[19788] <= 3'b110;
      // memory_array[19789] <= 3'b000;
      // memory_array[19790] <= 3'b000;
      // memory_array[19791] <= 3'b101;
      // memory_array[19792] <= 3'b101;
      // memory_array[19793] <= 3'b101;
      // memory_array[19794] <= 3'b000;
      // memory_array[19795] <= 3'b101;
      // memory_array[19796] <= 3'b101;
      // memory_array[19797] <= 3'b110;
      // memory_array[19798] <= 3'b101;
      // memory_array[19799] <= 3'b101;
      // memory_array[19800] <= 3'b101;
      // memory_array[19801] <= 3'b101;
      // memory_array[19802] <= 3'b101;
      // memory_array[19803] <= 3'b111;
      // memory_array[19804] <= 3'b111;
      // memory_array[19805] <= 3'b101;
      // memory_array[19806] <= 3'b101;
      // memory_array[19807] <= 3'b101;
      // memory_array[19808] <= 3'b101;
      // memory_array[19809] <= 3'b000;
      // memory_array[19810] <= 3'b000;
      // memory_array[19811] <= 3'b110;
      // memory_array[19812] <= 3'b000;
      // memory_array[19813] <= 3'b110;
      // memory_array[19814] <= 3'b110;
      // memory_array[19815] <= 3'b000;
      // memory_array[19816] <= 3'b110;
      // memory_array[19817] <= 3'b111;
      // memory_array[19818] <= 3'b110;
      // memory_array[19819] <= 3'b110;
      // memory_array[19820] <= 3'b111;
      // memory_array[19821] <= 3'b000;
      // memory_array[19822] <= 3'b110;
      // memory_array[19823] <= 3'b000;
      // memory_array[19824] <= 3'b111;
      // memory_array[19825] <= 3'b111;
      // memory_array[19826] <= 3'b111;
      // memory_array[19827] <= 3'b000;
      // memory_array[19828] <= 3'b110;
      // memory_array[19829] <= 3'b110;
      // memory_array[19830] <= 3'b111;
      // memory_array[19831] <= 3'b111;
      // memory_array[19832] <= 3'b000;
      // memory_array[19833] <= 3'b111;
      // memory_array[19834] <= 3'b111;
      // memory_array[19835] <= 3'b111;
      // memory_array[19836] <= 3'b000;
      // memory_array[19837] <= 3'b111;
      // memory_array[19838] <= 3'b111;
      // memory_array[19839] <= 3'b111;
      // memory_array[19840] <= 3'b111;
      // memory_array[19841] <= 3'b000;
      // memory_array[19842] <= 3'b000;
      // memory_array[19843] <= 3'b110;
      // memory_array[19844] <= 3'b111;
      // memory_array[19845] <= 3'b111;
      // memory_array[19846] <= 3'b111;
      // memory_array[19847] <= 3'b111;
      // memory_array[19848] <= 3'b111;
      // memory_array[19849] <= 3'b000;
      // memory_array[19850] <= 3'b000;
      // memory_array[19851] <= 3'b111;
      // memory_array[19852] <= 3'b111;
      // memory_array[19853] <= 3'b111;
      // memory_array[19854] <= 3'b111;
      // memory_array[19855] <= 3'b000;
      // memory_array[19856] <= 3'b000;
      // memory_array[19857] <= 3'b111;
      // memory_array[19858] <= 3'b111;
      // memory_array[19859] <= 3'b111;
      // memory_array[19860] <= 3'b111;
      // memory_array[19861] <= 3'b000;
      // memory_array[19862] <= 3'b000;
      // memory_array[19863] <= 3'b101;
      // memory_array[19864] <= 3'b101;
      // memory_array[19865] <= 3'b000;
      // memory_array[19866] <= 3'b000;
      // memory_array[19867] <= 3'b111;
      // memory_array[19868] <= 3'b111;
      // memory_array[19869] <= 3'b111;
      // memory_array[19870] <= 3'b111;
      // memory_array[19871] <= 3'b000;
      // memory_array[19872] <= 3'b111;
      // memory_array[19873] <= 3'b111;
      // memory_array[19874] <= 3'b111;
      // memory_array[19875] <= 3'b111;
      // memory_array[19876] <= 3'b000;
      // memory_array[19877] <= 3'b000;
      // memory_array[19878] <= 3'b000;
      // memory_array[19879] <= 3'b000;
      // memory_array[19880] <= 3'b000;
      // memory_array[19881] <= 3'b000;
      // memory_array[19882] <= 3'b111;
      // memory_array[19883] <= 3'b111;
      // memory_array[19884] <= 3'b111;
      // memory_array[19885] <= 3'b111;
      // memory_array[19886] <= 3'b000;
      // memory_array[19887] <= 3'b000;
      // memory_array[19888] <= 3'b101;
      // memory_array[19889] <= 3'b101;
      // memory_array[19890] <= 3'b000;
      // memory_array[19891] <= 3'b000;
      // memory_array[19892] <= 3'b000;
      // memory_array[19893] <= 3'b101;
      // memory_array[19894] <= 3'b000;
      // memory_array[19895] <= 3'b111;
      // memory_array[19896] <= 3'b111;
      // memory_array[19897] <= 3'b111;
      // memory_array[19898] <= 3'b111;
      // memory_array[19899] <= 3'b000;
      // memory_array[19900] <= 3'b000;
      // memory_array[19901] <= 3'b111;
      // memory_array[19902] <= 3'b111;
      // memory_array[19903] <= 3'b111;
      // memory_array[19904] <= 3'b000;
      // memory_array[19905] <= 3'b000;
      // memory_array[19906] <= 3'b000;
      // memory_array[19907] <= 3'b000;
      // memory_array[19908] <= 3'b111;
      // memory_array[19909] <= 3'b111;
      // memory_array[19910] <= 3'b111;
      // memory_array[19911] <= 3'b111;
      // memory_array[19912] <= 3'b111;
      // memory_array[19913] <= 3'b111;
      // memory_array[19914] <= 3'b111;
      // memory_array[19915] <= 3'b111;
      // memory_array[19916] <= 3'b000;
      // memory_array[19917] <= 3'b000;
      // memory_array[19918] <= 3'b101;
      // memory_array[19919] <= 3'b101;
      // memory_array[19920] <= 3'b101;
      // memory_array[19921] <= 3'b111;
      // memory_array[19922] <= 3'b111;
      // memory_array[19923] <= 3'b111;
      // memory_array[19924] <= 3'b111;
      // memory_array[19925] <= 3'b111;
      // memory_array[19926] <= 3'b000;
      // memory_array[19927] <= 3'b000;
      // memory_array[19928] <= 3'b101;
      // memory_array[19929] <= 3'b000;
      // memory_array[19930] <= 3'b000;
      // memory_array[19931] <= 3'b000;
      // memory_array[19932] <= 3'b000;
      // memory_array[19933] <= 3'b101;
      // memory_array[19934] <= 3'b000;
      // memory_array[19935] <= 3'b111;
      // memory_array[19936] <= 3'b111;
      // memory_array[19937] <= 3'b111;
      // memory_array[19938] <= 3'b111;
      // memory_array[19939] <= 3'b111;
      // memory_array[19940] <= 3'b111;
      // memory_array[19941] <= 3'b111;
      // memory_array[19942] <= 3'b000;
      // memory_array[19943] <= 3'b000;
      // memory_array[19944] <= 3'b101;
      // memory_array[19945] <= 3'b000;
      // memory_array[19946] <= 3'b000;
      // memory_array[19947] <= 3'b000;
      // memory_array[19948] <= 3'b101;
      // memory_array[19949] <= 3'b111;
      // memory_array[19950] <= 3'b111;
      // memory_array[19951] <= 3'b000;
      // memory_array[19952] <= 3'b000;
      // memory_array[19953] <= 3'b111;
      // memory_array[19954] <= 3'b111;
      // memory_array[19955] <= 3'b111;
      // memory_array[19956] <= 3'b111;
      // memory_array[19957] <= 3'b111;
      // memory_array[19958] <= 3'b111;
      // memory_array[19959] <= 3'b110;
      // memory_array[19960] <= 3'b000;
      // memory_array[19961] <= 3'b000;
      // memory_array[19962] <= 3'b111;
      // memory_array[19963] <= 3'b111;
      // memory_array[19964] <= 3'b111;
      // memory_array[19965] <= 3'b111;
      // memory_array[19966] <= 3'b110;
      // memory_array[19967] <= 3'b111;
      // memory_array[19968] <= 3'b110;
      // memory_array[19969] <= 3'b110;
      // memory_array[19970] <= 3'b110;
      // memory_array[19971] <= 3'b111;
      // memory_array[19972] <= 3'b111;
      // memory_array[19973] <= 3'b111;
      // memory_array[19974] <= 3'b111;
      // memory_array[19975] <= 3'b111;
      // memory_array[19976] <= 3'b111;
      // memory_array[19977] <= 3'b111;
      // memory_array[19978] <= 3'b111;
      // memory_array[19979] <= 3'b110;
      // memory_array[19980] <= 3'b110;
      // memory_array[19981] <= 3'b110;
      // memory_array[19982] <= 3'b110;
      // memory_array[19983] <= 3'b110;
      // memory_array[19984] <= 3'b110;
      // memory_array[19985] <= 3'b000;
      // memory_array[19986] <= 3'b000;
      // memory_array[19987] <= 3'b000;
      // memory_array[19988] <= 3'b110;
      // memory_array[19989] <= 3'b000;
      // memory_array[19990] <= 3'b000;
      // memory_array[19991] <= 3'b101;
      // memory_array[19992] <= 3'b101;
      // memory_array[19993] <= 3'b101;
      // memory_array[19994] <= 3'b101;
      // memory_array[19995] <= 3'b111;
      // memory_array[19996] <= 3'b111;
      // memory_array[19997] <= 3'b101;
      // memory_array[19998] <= 3'b101;
      // memory_array[19999] <= 3'b101;
      // memory_array[20000] <= 3'b101;
      // memory_array[20001] <= 3'b101;
      // memory_array[20002] <= 3'b101;
      // memory_array[20003] <= 3'b101;
      // memory_array[20004] <= 3'b101;
      // memory_array[20005] <= 3'b101;
      // memory_array[20006] <= 3'b101;
      // memory_array[20007] <= 3'b101;
      // memory_array[20008] <= 3'b101;
      // memory_array[20009] <= 3'b000;
      // memory_array[20010] <= 3'b000;
      // memory_array[20011] <= 3'b110;
      // memory_array[20012] <= 3'b110;
      // memory_array[20013] <= 3'b000;
      // memory_array[20014] <= 3'b000;
      // memory_array[20015] <= 3'b110;
      // memory_array[20016] <= 3'b110;
      // memory_array[20017] <= 3'b110;
      // memory_array[20018] <= 3'b111;
      // memory_array[20019] <= 3'b111;
      // memory_array[20020] <= 3'b110;
      // memory_array[20021] <= 3'b000;
      // memory_array[20022] <= 3'b110;
      // memory_array[20023] <= 3'b000;
      // memory_array[20024] <= 3'b111;
      // memory_array[20025] <= 3'b111;
      // memory_array[20026] <= 3'b111;
      // memory_array[20027] <= 3'b000;
      // memory_array[20028] <= 3'b111;
      // memory_array[20029] <= 3'b111;
      // memory_array[20030] <= 3'b110;
      // memory_array[20031] <= 3'b110;
      // memory_array[20032] <= 3'b000;
      // memory_array[20033] <= 3'b111;
      // memory_array[20034] <= 3'b111;
      // memory_array[20035] <= 3'b111;
      // memory_array[20036] <= 3'b110;
      // memory_array[20037] <= 3'b111;
      // memory_array[20038] <= 3'b111;
      // memory_array[20039] <= 3'b111;
      // memory_array[20040] <= 3'b111;
      // memory_array[20041] <= 3'b000;
      // memory_array[20042] <= 3'b000;
      // memory_array[20043] <= 3'b000;
      // memory_array[20044] <= 3'b111;
      // memory_array[20045] <= 3'b111;
      // memory_array[20046] <= 3'b111;
      // memory_array[20047] <= 3'b111;
      // memory_array[20048] <= 3'b000;
      // memory_array[20049] <= 3'b000;
      // memory_array[20050] <= 3'b000;
      // memory_array[20051] <= 3'b111;
      // memory_array[20052] <= 3'b111;
      // memory_array[20053] <= 3'b111;
      // memory_array[20054] <= 3'b111;
      // memory_array[20055] <= 3'b000;
      // memory_array[20056] <= 3'b000;
      // memory_array[20057] <= 3'b111;
      // memory_array[20058] <= 3'b111;
      // memory_array[20059] <= 3'b111;
      // memory_array[20060] <= 3'b111;
      // memory_array[20061] <= 3'b000;
      // memory_array[20062] <= 3'b101;
      // memory_array[20063] <= 3'b000;
      // memory_array[20064] <= 3'b000;
      // memory_array[20065] <= 3'b101;
      // memory_array[20066] <= 3'b000;
      // memory_array[20067] <= 3'b111;
      // memory_array[20068] <= 3'b111;
      // memory_array[20069] <= 3'b111;
      // memory_array[20070] <= 3'b111;
      // memory_array[20071] <= 3'b000;
      // memory_array[20072] <= 3'b111;
      // memory_array[20073] <= 3'b111;
      // memory_array[20074] <= 3'b111;
      // memory_array[20075] <= 3'b111;
      // memory_array[20076] <= 3'b000;
      // memory_array[20077] <= 3'b000;
      // memory_array[20078] <= 3'b000;
      // memory_array[20079] <= 3'b000;
      // memory_array[20080] <= 3'b000;
      // memory_array[20081] <= 3'b000;
      // memory_array[20082] <= 3'b111;
      // memory_array[20083] <= 3'b111;
      // memory_array[20084] <= 3'b111;
      // memory_array[20085] <= 3'b111;
      // memory_array[20086] <= 3'b111;
      // memory_array[20087] <= 3'b101;
      // memory_array[20088] <= 3'b000;
      // memory_array[20089] <= 3'b000;
      // memory_array[20090] <= 3'b101;
      // memory_array[20091] <= 3'b101;
      // memory_array[20092] <= 3'b101;
      // memory_array[20093] <= 3'b000;
      // memory_array[20094] <= 3'b000;
      // memory_array[20095] <= 3'b000;
      // memory_array[20096] <= 3'b111;
      // memory_array[20097] <= 3'b111;
      // memory_array[20098] <= 3'b111;
      // memory_array[20099] <= 3'b110;
      // memory_array[20100] <= 3'b110;
      // memory_array[20101] <= 3'b111;
      // memory_array[20102] <= 3'b111;
      // memory_array[20103] <= 3'b111;
      // memory_array[20104] <= 3'b000;
      // memory_array[20105] <= 3'b000;
      // memory_array[20106] <= 3'b101;
      // memory_array[20107] <= 3'b000;
      // memory_array[20108] <= 3'b111;
      // memory_array[20109] <= 3'b111;
      // memory_array[20110] <= 3'b111;
      // memory_array[20111] <= 3'b111;
      // memory_array[20112] <= 3'b000;
      // memory_array[20113] <= 3'b000;
      // memory_array[20114] <= 3'b111;
      // memory_array[20115] <= 3'b000;
      // memory_array[20116] <= 3'b101;
      // memory_array[20117] <= 3'b101;
      // memory_array[20118] <= 3'b101;
      // memory_array[20119] <= 3'b101;
      // memory_array[20120] <= 3'b000;
      // memory_array[20121] <= 3'b111;
      // memory_array[20122] <= 3'b111;
      // memory_array[20123] <= 3'b111;
      // memory_array[20124] <= 3'b111;
      // memory_array[20125] <= 3'b111;
      // memory_array[20126] <= 3'b101;
      // memory_array[20127] <= 3'b101;
      // memory_array[20128] <= 3'b000;
      // memory_array[20129] <= 3'b000;
      // memory_array[20130] <= 3'b000;
      // memory_array[20131] <= 3'b000;
      // memory_array[20132] <= 3'b000;
      // memory_array[20133] <= 3'b000;
      // memory_array[20134] <= 3'b000;
      // memory_array[20135] <= 3'b111;
      // memory_array[20136] <= 3'b111;
      // memory_array[20137] <= 3'b111;
      // memory_array[20138] <= 3'b111;
      // memory_array[20139] <= 3'b111;
      // memory_array[20140] <= 3'b111;
      // memory_array[20141] <= 3'b111;
      // memory_array[20142] <= 3'b111;
      // memory_array[20143] <= 3'b000;
      // memory_array[20144] <= 3'b000;
      // memory_array[20145] <= 3'b101;
      // memory_array[20146] <= 3'b101;
      // memory_array[20147] <= 3'b101;
      // memory_array[20148] <= 3'b000;
      // memory_array[20149] <= 3'b111;
      // memory_array[20150] <= 3'b111;
      // memory_array[20151] <= 3'b111;
      // memory_array[20152] <= 3'b000;
      // memory_array[20153] <= 3'b000;
      // memory_array[20154] <= 3'b111;
      // memory_array[20155] <= 3'b111;
      // memory_array[20156] <= 3'b111;
      // memory_array[20157] <= 3'b111;
      // memory_array[20158] <= 3'b111;
      // memory_array[20159] <= 3'b000;
      // memory_array[20160] <= 3'b110;
      // memory_array[20161] <= 3'b000;
      // memory_array[20162] <= 3'b111;
      // memory_array[20163] <= 3'b111;
      // memory_array[20164] <= 3'b111;
      // memory_array[20165] <= 3'b111;
      // memory_array[20166] <= 3'b110;
      // memory_array[20167] <= 3'b110;
      // memory_array[20168] <= 3'b110;
      // memory_array[20169] <= 3'b110;
      // memory_array[20170] <= 3'b000;
      // memory_array[20171] <= 3'b111;
      // memory_array[20172] <= 3'b111;
      // memory_array[20173] <= 3'b111;
      // memory_array[20174] <= 3'b000;
      // memory_array[20175] <= 3'b111;
      // memory_array[20176] <= 3'b111;
      // memory_array[20177] <= 3'b111;
      // memory_array[20178] <= 3'b111;
      // memory_array[20179] <= 3'b110;
      // memory_array[20180] <= 3'b110;
      // memory_array[20181] <= 3'b110;
      // memory_array[20182] <= 3'b110;
      // memory_array[20183] <= 3'b000;
      // memory_array[20184] <= 3'b110;
      // memory_array[20185] <= 3'b110;
      // memory_array[20186] <= 3'b110;
      // memory_array[20187] <= 3'b110;
      // memory_array[20188] <= 3'b000;
      // memory_array[20189] <= 3'b000;
      // memory_array[20190] <= 3'b000;
      // memory_array[20191] <= 3'b101;
      // memory_array[20192] <= 3'b101;
      // memory_array[20193] <= 3'b101;
      // memory_array[20194] <= 3'b101;
      // memory_array[20195] <= 3'b101;
      // memory_array[20196] <= 3'b101;
      // memory_array[20197] <= 3'b101;
      // memory_array[20198] <= 3'b101;
      // memory_array[20199] <= 3'b101;
      // memory_array[20200] <= 3'b101;
      // memory_array[20201] <= 3'b101;
      // memory_array[20202] <= 3'b101;
      // memory_array[20203] <= 3'b101;
      // memory_array[20204] <= 3'b101;
      // memory_array[20205] <= 3'b101;
      // memory_array[20206] <= 3'b101;
      // memory_array[20207] <= 3'b101;
      // memory_array[20208] <= 3'b101;
      // memory_array[20209] <= 3'b000;
      // memory_array[20210] <= 3'b000;
      // memory_array[20211] <= 3'b110;
      // memory_array[20212] <= 3'b110;
      // memory_array[20213] <= 3'b000;
      // memory_array[20214] <= 3'b000;
      // memory_array[20215] <= 3'b110;
      // memory_array[20216] <= 3'b110;
      // memory_array[20217] <= 3'b110;
      // memory_array[20218] <= 3'b111;
      // memory_array[20219] <= 3'b111;
      // memory_array[20220] <= 3'b110;
      // memory_array[20221] <= 3'b000;
      // memory_array[20222] <= 3'b110;
      // memory_array[20223] <= 3'b000;
      // memory_array[20224] <= 3'b111;
      // memory_array[20225] <= 3'b111;
      // memory_array[20226] <= 3'b111;
      // memory_array[20227] <= 3'b000;
      // memory_array[20228] <= 3'b111;
      // memory_array[20229] <= 3'b111;
      // memory_array[20230] <= 3'b110;
      // memory_array[20231] <= 3'b110;
      // memory_array[20232] <= 3'b111;
      // memory_array[20233] <= 3'b111;
      // memory_array[20234] <= 3'b111;
      // memory_array[20235] <= 3'b000;
      // memory_array[20236] <= 3'b110;
      // memory_array[20237] <= 3'b111;
      // memory_array[20238] <= 3'b111;
      // memory_array[20239] <= 3'b111;
      // memory_array[20240] <= 3'b111;
      // memory_array[20241] <= 3'b111;
      // memory_array[20242] <= 3'b111;
      // memory_array[20243] <= 3'b111;
      // memory_array[20244] <= 3'b111;
      // memory_array[20245] <= 3'b111;
      // memory_array[20246] <= 3'b111;
      // memory_array[20247] <= 3'b111;
      // memory_array[20248] <= 3'b111;
      // memory_array[20249] <= 3'b101;
      // memory_array[20250] <= 3'b000;
      // memory_array[20251] <= 3'b111;
      // memory_array[20252] <= 3'b111;
      // memory_array[20253] <= 3'b111;
      // memory_array[20254] <= 3'b111;
      // memory_array[20255] <= 3'b000;
      // memory_array[20256] <= 3'b000;
      // memory_array[20257] <= 3'b111;
      // memory_array[20258] <= 3'b111;
      // memory_array[20259] <= 3'b111;
      // memory_array[20260] <= 3'b111;
      // memory_array[20261] <= 3'b000;
      // memory_array[20262] <= 3'b000;
      // memory_array[20263] <= 3'b000;
      // memory_array[20264] <= 3'b000;
      // memory_array[20265] <= 3'b101;
      // memory_array[20266] <= 3'b000;
      // memory_array[20267] <= 3'b111;
      // memory_array[20268] <= 3'b111;
      // memory_array[20269] <= 3'b111;
      // memory_array[20270] <= 3'b111;
      // memory_array[20271] <= 3'b000;
      // memory_array[20272] <= 3'b111;
      // memory_array[20273] <= 3'b111;
      // memory_array[20274] <= 3'b111;
      // memory_array[20275] <= 3'b111;
      // memory_array[20276] <= 3'b000;
      // memory_array[20277] <= 3'b000;
      // memory_array[20278] <= 3'b000;
      // memory_array[20279] <= 3'b000;
      // memory_array[20280] <= 3'b000;
      // memory_array[20281] <= 3'b000;
      // memory_array[20282] <= 3'b000;
      // memory_array[20283] <= 3'b111;
      // memory_array[20284] <= 3'b111;
      // memory_array[20285] <= 3'b111;
      // memory_array[20286] <= 3'b111;
      // memory_array[20287] <= 3'b101;
      // memory_array[20288] <= 3'b000;
      // memory_array[20289] <= 3'b000;
      // memory_array[20290] <= 3'b101;
      // memory_array[20291] <= 3'b000;
      // memory_array[20292] <= 3'b111;
      // memory_array[20293] <= 3'b111;
      // memory_array[20294] <= 3'b111;
      // memory_array[20295] <= 3'b111;
      // memory_array[20296] <= 3'b000;
      // memory_array[20297] <= 3'b101;
      // memory_array[20298] <= 3'b000;
      // memory_array[20299] <= 3'b000;
      // memory_array[20300] <= 3'b110;
      // memory_array[20301] <= 3'b111;
      // memory_array[20302] <= 3'b111;
      // memory_array[20303] <= 3'b111;
      // memory_array[20304] <= 3'b000;
      // memory_array[20305] <= 3'b101;
      // memory_array[20306] <= 3'b000;
      // memory_array[20307] <= 3'b000;
      // memory_array[20308] <= 3'b111;
      // memory_array[20309] <= 3'b111;
      // memory_array[20310] <= 3'b111;
      // memory_array[20311] <= 3'b111;
      // memory_array[20312] <= 3'b101;
      // memory_array[20313] <= 3'b101;
      // memory_array[20314] <= 3'b000;
      // memory_array[20315] <= 3'b101;
      // memory_array[20316] <= 3'b000;
      // memory_array[20317] <= 3'b101;
      // memory_array[20318] <= 3'b000;
      // memory_array[20319] <= 3'b000;
      // memory_array[20320] <= 3'b000;
      // memory_array[20321] <= 3'b000;
      // memory_array[20322] <= 3'b111;
      // memory_array[20323] <= 3'b111;
      // memory_array[20324] <= 3'b111;
      // memory_array[20325] <= 3'b111;
      // memory_array[20326] <= 3'b000;
      // memory_array[20327] <= 3'b000;
      // memory_array[20328] <= 3'b000;
      // memory_array[20329] <= 3'b000;
      // memory_array[20330] <= 3'b111;
      // memory_array[20331] <= 3'b111;
      // memory_array[20332] <= 3'b111;
      // memory_array[20333] <= 3'b111;
      // memory_array[20334] <= 3'b111;
      // memory_array[20335] <= 3'b111;
      // memory_array[20336] <= 3'b111;
      // memory_array[20337] <= 3'b111;
      // memory_array[20338] <= 3'b111;
      // memory_array[20339] <= 3'b111;
      // memory_array[20340] <= 3'b111;
      // memory_array[20341] <= 3'b111;
      // memory_array[20342] <= 3'b111;
      // memory_array[20343] <= 3'b111;
      // memory_array[20344] <= 3'b000;
      // memory_array[20345] <= 3'b000;
      // memory_array[20346] <= 3'b101;
      // memory_array[20347] <= 3'b101;
      // memory_array[20348] <= 3'b000;
      // memory_array[20349] <= 3'b111;
      // memory_array[20350] <= 3'b111;
      // memory_array[20351] <= 3'b111;
      // memory_array[20352] <= 3'b000;
      // memory_array[20353] <= 3'b111;
      // memory_array[20354] <= 3'b111;
      // memory_array[20355] <= 3'b111;
      // memory_array[20356] <= 3'b111;
      // memory_array[20357] <= 3'b111;
      // memory_array[20358] <= 3'b111;
      // memory_array[20359] <= 3'b111;
      // memory_array[20360] <= 3'b000;
      // memory_array[20361] <= 3'b000;
      // memory_array[20362] <= 3'b111;
      // memory_array[20363] <= 3'b111;
      // memory_array[20364] <= 3'b111;
      // memory_array[20365] <= 3'b111;
      // memory_array[20366] <= 3'b110;
      // memory_array[20367] <= 3'b110;
      // memory_array[20368] <= 3'b110;
      // memory_array[20369] <= 3'b111;
      // memory_array[20370] <= 3'b111;
      // memory_array[20371] <= 3'b111;
      // memory_array[20372] <= 3'b000;
      // memory_array[20373] <= 3'b110;
      // memory_array[20374] <= 3'b000;
      // memory_array[20375] <= 3'b111;
      // memory_array[20376] <= 3'b111;
      // memory_array[20377] <= 3'b111;
      // memory_array[20378] <= 3'b111;
      // memory_array[20379] <= 3'b110;
      // memory_array[20380] <= 3'b110;
      // memory_array[20381] <= 3'b110;
      // memory_array[20382] <= 3'b110;
      // memory_array[20383] <= 3'b000;
      // memory_array[20384] <= 3'b110;
      // memory_array[20385] <= 3'b110;
      // memory_array[20386] <= 3'b110;
      // memory_array[20387] <= 3'b110;
      // memory_array[20388] <= 3'b000;
      // memory_array[20389] <= 3'b000;
      // memory_array[20390] <= 3'b000;
      // memory_array[20391] <= 3'b101;
      // memory_array[20392] <= 3'b101;
      // memory_array[20393] <= 3'b101;
      // memory_array[20394] <= 3'b101;
      // memory_array[20395] <= 3'b101;
      // memory_array[20396] <= 3'b101;
      // memory_array[20397] <= 3'b101;
      // memory_array[20398] <= 3'b101;
      // memory_array[20399] <= 3'b101;
      // memory_array[20400] <= 3'b101;
      // memory_array[20401] <= 3'b101;
      // memory_array[20402] <= 3'b101;
      // memory_array[20403] <= 3'b111;
      // memory_array[20404] <= 3'b111;
      // memory_array[20405] <= 3'b101;
      // memory_array[20406] <= 3'b101;
      // memory_array[20407] <= 3'b101;
      // memory_array[20408] <= 3'b101;
      // memory_array[20409] <= 3'b000;
      // memory_array[20410] <= 3'b000;
      // memory_array[20411] <= 3'b110;
      // memory_array[20412] <= 3'b000;
      // memory_array[20413] <= 3'b110;
      // memory_array[20414] <= 3'b110;
      // memory_array[20415] <= 3'b000;
      // memory_array[20416] <= 3'b110;
      // memory_array[20417] <= 3'b111;
      // memory_array[20418] <= 3'b110;
      // memory_array[20419] <= 3'b110;
      // memory_array[20420] <= 3'b111;
      // memory_array[20421] <= 3'b000;
      // memory_array[20422] <= 3'b110;
      // memory_array[20423] <= 3'b000;
      // memory_array[20424] <= 3'b111;
      // memory_array[20425] <= 3'b111;
      // memory_array[20426] <= 3'b111;
      // memory_array[20427] <= 3'b000;
      // memory_array[20428] <= 3'b110;
      // memory_array[20429] <= 3'b110;
      // memory_array[20430] <= 3'b111;
      // memory_array[20431] <= 3'b000;
      // memory_array[20432] <= 3'b111;
      // memory_array[20433] <= 3'b111;
      // memory_array[20434] <= 3'b111;
      // memory_array[20435] <= 3'b000;
      // memory_array[20436] <= 3'b110;
      // memory_array[20437] <= 3'b111;
      // memory_array[20438] <= 3'b111;
      // memory_array[20439] <= 3'b111;
      // memory_array[20440] <= 3'b111;
      // memory_array[20441] <= 3'b111;
      // memory_array[20442] <= 3'b111;
      // memory_array[20443] <= 3'b111;
      // memory_array[20444] <= 3'b111;
      // memory_array[20445] <= 3'b111;
      // memory_array[20446] <= 3'b000;
      // memory_array[20447] <= 3'b111;
      // memory_array[20448] <= 3'b111;
      // memory_array[20449] <= 3'b101;
      // memory_array[20450] <= 3'b000;
      // memory_array[20451] <= 3'b111;
      // memory_array[20452] <= 3'b111;
      // memory_array[20453] <= 3'b111;
      // memory_array[20454] <= 3'b111;
      // memory_array[20455] <= 3'b000;
      // memory_array[20456] <= 3'b000;
      // memory_array[20457] <= 3'b111;
      // memory_array[20458] <= 3'b111;
      // memory_array[20459] <= 3'b111;
      // memory_array[20460] <= 3'b111;
      // memory_array[20461] <= 3'b000;
      // memory_array[20462] <= 3'b000;
      // memory_array[20463] <= 3'b101;
      // memory_array[20464] <= 3'b101;
      // memory_array[20465] <= 3'b000;
      // memory_array[20466] <= 3'b000;
      // memory_array[20467] <= 3'b111;
      // memory_array[20468] <= 3'b111;
      // memory_array[20469] <= 3'b111;
      // memory_array[20470] <= 3'b111;
      // memory_array[20471] <= 3'b000;
      // memory_array[20472] <= 3'b000;
      // memory_array[20473] <= 3'b111;
      // memory_array[20474] <= 3'b111;
      // memory_array[20475] <= 3'b111;
      // memory_array[20476] <= 3'b111;
      // memory_array[20477] <= 3'b000;
      // memory_array[20478] <= 3'b000;
      // memory_array[20479] <= 3'b000;
      // memory_array[20480] <= 3'b000;
      // memory_array[20481] <= 3'b000;
      // memory_array[20482] <= 3'b000;
      // memory_array[20483] <= 3'b111;
      // memory_array[20484] <= 3'b111;
      // memory_array[20485] <= 3'b111;
      // memory_array[20486] <= 3'b111;
      // memory_array[20487] <= 3'b000;
      // memory_array[20488] <= 3'b101;
      // memory_array[20489] <= 3'b101;
      // memory_array[20490] <= 3'b000;
      // memory_array[20491] <= 3'b000;
      // memory_array[20492] <= 3'b111;
      // memory_array[20493] <= 3'b111;
      // memory_array[20494] <= 3'b111;
      // memory_array[20495] <= 3'b111;
      // memory_array[20496] <= 3'b000;
      // memory_array[20497] <= 3'b000;
      // memory_array[20498] <= 3'b101;
      // memory_array[20499] <= 3'b000;
      // memory_array[20500] <= 3'b000;
      // memory_array[20501] <= 3'b111;
      // memory_array[20502] <= 3'b111;
      // memory_array[20503] <= 3'b111;
      // memory_array[20504] <= 3'b000;
      // memory_array[20505] <= 3'b000;
      // memory_array[20506] <= 3'b000;
      // memory_array[20507] <= 3'b000;
      // memory_array[20508] <= 3'b111;
      // memory_array[20509] <= 3'b111;
      // memory_array[20510] <= 3'b111;
      // memory_array[20511] <= 3'b111;
      // memory_array[20512] <= 3'b101;
      // memory_array[20513] <= 3'b101;
      // memory_array[20514] <= 3'b101;
      // memory_array[20515] <= 3'b101;
      // memory_array[20516] <= 3'b000;
      // memory_array[20517] <= 3'b000;
      // memory_array[20518] <= 3'b000;
      // memory_array[20519] <= 3'b000;
      // memory_array[20520] <= 3'b000;
      // memory_array[20521] <= 3'b000;
      // memory_array[20522] <= 3'b111;
      // memory_array[20523] <= 3'b111;
      // memory_array[20524] <= 3'b111;
      // memory_array[20525] <= 3'b111;
      // memory_array[20526] <= 3'b000;
      // memory_array[20527] <= 3'b000;
      // memory_array[20528] <= 3'b000;
      // memory_array[20529] <= 3'b000;
      // memory_array[20530] <= 3'b000;
      // memory_array[20531] <= 3'b111;
      // memory_array[20532] <= 3'b111;
      // memory_array[20533] <= 3'b111;
      // memory_array[20534] <= 3'b111;
      // memory_array[20535] <= 3'b111;
      // memory_array[20536] <= 3'b111;
      // memory_array[20537] <= 3'b111;
      // memory_array[20538] <= 3'b111;
      // memory_array[20539] <= 3'b000;
      // memory_array[20540] <= 3'b111;
      // memory_array[20541] <= 3'b111;
      // memory_array[20542] <= 3'b111;
      // memory_array[20543] <= 3'b111;
      // memory_array[20544] <= 3'b000;
      // memory_array[20545] <= 3'b000;
      // memory_array[20546] <= 3'b000;
      // memory_array[20547] <= 3'b000;
      // memory_array[20548] <= 3'b111;
      // memory_array[20549] <= 3'b111;
      // memory_array[20550] <= 3'b111;
      // memory_array[20551] <= 3'b111;
      // memory_array[20552] <= 3'b000;
      // memory_array[20553] <= 3'b111;
      // memory_array[20554] <= 3'b000;
      // memory_array[20555] <= 3'b111;
      // memory_array[20556] <= 3'b111;
      // memory_array[20557] <= 3'b111;
      // memory_array[20558] <= 3'b111;
      // memory_array[20559] <= 3'b111;
      // memory_array[20560] <= 3'b000;
      // memory_array[20561] <= 3'b000;
      // memory_array[20562] <= 3'b111;
      // memory_array[20563] <= 3'b111;
      // memory_array[20564] <= 3'b111;
      // memory_array[20565] <= 3'b111;
      // memory_array[20566] <= 3'b110;
      // memory_array[20567] <= 3'b111;
      // memory_array[20568] <= 3'b000;
      // memory_array[20569] <= 3'b111;
      // memory_array[20570] <= 3'b111;
      // memory_array[20571] <= 3'b111;
      // memory_array[20572] <= 3'b000;
      // memory_array[20573] <= 3'b110;
      // memory_array[20574] <= 3'b000;
      // memory_array[20575] <= 3'b111;
      // memory_array[20576] <= 3'b111;
      // memory_array[20577] <= 3'b111;
      // memory_array[20578] <= 3'b111;
      // memory_array[20579] <= 3'b110;
      // memory_array[20580] <= 3'b110;
      // memory_array[20581] <= 3'b110;
      // memory_array[20582] <= 3'b110;
      // memory_array[20583] <= 3'b110;
      // memory_array[20584] <= 3'b110;
      // memory_array[20585] <= 3'b000;
      // memory_array[20586] <= 3'b000;
      // memory_array[20587] <= 3'b000;
      // memory_array[20588] <= 3'b110;
      // memory_array[20589] <= 3'b000;
      // memory_array[20590] <= 3'b000;
      // memory_array[20591] <= 3'b101;
      // memory_array[20592] <= 3'b101;
      // memory_array[20593] <= 3'b101;
      // memory_array[20594] <= 3'b101;
      // memory_array[20595] <= 3'b111;
      // memory_array[20596] <= 3'b111;
      // memory_array[20597] <= 3'b101;
      // memory_array[20598] <= 3'b101;
      // memory_array[20599] <= 3'b101;
      // memory_array[20600] <= 3'b101;
      // memory_array[20601] <= 3'b101;
      // memory_array[20602] <= 3'b110;
      // memory_array[20603] <= 3'b101;
      // memory_array[20604] <= 3'b101;
      // memory_array[20605] <= 3'b110;
      // memory_array[20606] <= 3'b101;
      // memory_array[20607] <= 3'b101;
      // memory_array[20608] <= 3'b101;
      // memory_array[20609] <= 3'b000;
      // memory_array[20610] <= 3'b000;
      // memory_array[20611] <= 3'b110;
      // memory_array[20612] <= 3'b110;
      // memory_array[20613] <= 3'b000;
      // memory_array[20614] <= 3'b000;
      // memory_array[20615] <= 3'b000;
      // memory_array[20616] <= 3'b110;
      // memory_array[20617] <= 3'b110;
      // memory_array[20618] <= 3'b110;
      // memory_array[20619] <= 3'b110;
      // memory_array[20620] <= 3'b110;
      // memory_array[20621] <= 3'b000;
      // memory_array[20622] <= 3'b110;
      // memory_array[20623] <= 3'b000;
      // memory_array[20624] <= 3'b111;
      // memory_array[20625] <= 3'b111;
      // memory_array[20626] <= 3'b111;
      // memory_array[20627] <= 3'b000;
      // memory_array[20628] <= 3'b111;
      // memory_array[20629] <= 3'b110;
      // memory_array[20630] <= 3'b110;
      // memory_array[20631] <= 3'b111;
      // memory_array[20632] <= 3'b111;
      // memory_array[20633] <= 3'b111;
      // memory_array[20634] <= 3'b000;
      // memory_array[20635] <= 3'b110;
      // memory_array[20636] <= 3'b110;
      // memory_array[20637] <= 3'b111;
      // memory_array[20638] <= 3'b111;
      // memory_array[20639] <= 3'b111;
      // memory_array[20640] <= 3'b111;
      // memory_array[20641] <= 3'b111;
      // memory_array[20642] <= 3'b111;
      // memory_array[20643] <= 3'b111;
      // memory_array[20644] <= 3'b000;
      // memory_array[20645] <= 3'b000;
      // memory_array[20646] <= 3'b111;
      // memory_array[20647] <= 3'b111;
      // memory_array[20648] <= 3'b111;
      // memory_array[20649] <= 3'b101;
      // memory_array[20650] <= 3'b000;
      // memory_array[20651] <= 3'b111;
      // memory_array[20652] <= 3'b111;
      // memory_array[20653] <= 3'b111;
      // memory_array[20654] <= 3'b111;
      // memory_array[20655] <= 3'b000;
      // memory_array[20656] <= 3'b101;
      // memory_array[20657] <= 3'b111;
      // memory_array[20658] <= 3'b111;
      // memory_array[20659] <= 3'b111;
      // memory_array[20660] <= 3'b111;
      // memory_array[20661] <= 3'b000;
      // memory_array[20662] <= 3'b101;
      // memory_array[20663] <= 3'b000;
      // memory_array[20664] <= 3'b000;
      // memory_array[20665] <= 3'b101;
      // memory_array[20666] <= 3'b101;
      // memory_array[20667] <= 3'b111;
      // memory_array[20668] <= 3'b111;
      // memory_array[20669] <= 3'b111;
      // memory_array[20670] <= 3'b111;
      // memory_array[20671] <= 3'b000;
      // memory_array[20672] <= 3'b000;
      // memory_array[20673] <= 3'b111;
      // memory_array[20674] <= 3'b111;
      // memory_array[20675] <= 3'b111;
      // memory_array[20676] <= 3'b111;
      // memory_array[20677] <= 3'b000;
      // memory_array[20678] <= 3'b000;
      // memory_array[20679] <= 3'b000;
      // memory_array[20680] <= 3'b000;
      // memory_array[20681] <= 3'b000;
      // memory_array[20682] <= 3'b000;
      // memory_array[20683] <= 3'b000;
      // memory_array[20684] <= 3'b111;
      // memory_array[20685] <= 3'b111;
      // memory_array[20686] <= 3'b111;
      // memory_array[20687] <= 3'b000;
      // memory_array[20688] <= 3'b000;
      // memory_array[20689] <= 3'b110;
      // memory_array[20690] <= 3'b101;
      // memory_array[20691] <= 3'b101;
      // memory_array[20692] <= 3'b111;
      // memory_array[20693] <= 3'b111;
      // memory_array[20694] <= 3'b111;
      // memory_array[20695] <= 3'b111;
      // memory_array[20696] <= 3'b000;
      // memory_array[20697] <= 3'b101;
      // memory_array[20698] <= 3'b000;
      // memory_array[20699] <= 3'b000;
      // memory_array[20700] <= 3'b110;
      // memory_array[20701] <= 3'b111;
      // memory_array[20702] <= 3'b111;
      // memory_array[20703] <= 3'b111;
      // memory_array[20704] <= 3'b000;
      // memory_array[20705] <= 3'b000;
      // memory_array[20706] <= 3'b101;
      // memory_array[20707] <= 3'b000;
      // memory_array[20708] <= 3'b111;
      // memory_array[20709] <= 3'b111;
      // memory_array[20710] <= 3'b111;
      // memory_array[20711] <= 3'b111;
      // memory_array[20712] <= 3'b101;
      // memory_array[20713] <= 3'b101;
      // memory_array[20714] <= 3'b101;
      // memory_array[20715] <= 3'b101;
      // memory_array[20716] <= 3'b000;
      // memory_array[20717] <= 3'b101;
      // memory_array[20718] <= 3'b000;
      // memory_array[20719] <= 3'b000;
      // memory_array[20720] <= 3'b000;
      // memory_array[20721] <= 3'b000;
      // memory_array[20722] <= 3'b111;
      // memory_array[20723] <= 3'b111;
      // memory_array[20724] <= 3'b111;
      // memory_array[20725] <= 3'b111;
      // memory_array[20726] <= 3'b111;
      // memory_array[20727] <= 3'b000;
      // memory_array[20728] <= 3'b000;
      // memory_array[20729] <= 3'b000;
      // memory_array[20730] <= 3'b000;
      // memory_array[20731] <= 3'b111;
      // memory_array[20732] <= 3'b111;
      // memory_array[20733] <= 3'b111;
      // memory_array[20734] <= 3'b000;
      // memory_array[20735] <= 3'b111;
      // memory_array[20736] <= 3'b111;
      // memory_array[20737] <= 3'b111;
      // memory_array[20738] <= 3'b111;
      // memory_array[20739] <= 3'b000;
      // memory_array[20740] <= 3'b000;
      // memory_array[20741] <= 3'b111;
      // memory_array[20742] <= 3'b111;
      // memory_array[20743] <= 3'b111;
      // memory_array[20744] <= 3'b000;
      // memory_array[20745] <= 3'b000;
      // memory_array[20746] <= 3'b000;
      // memory_array[20747] <= 3'b111;
      // memory_array[20748] <= 3'b111;
      // memory_array[20749] <= 3'b111;
      // memory_array[20750] <= 3'b111;
      // memory_array[20751] <= 3'b111;
      // memory_array[20752] <= 3'b111;
      // memory_array[20753] <= 3'b000;
      // memory_array[20754] <= 3'b111;
      // memory_array[20755] <= 3'b000;
      // memory_array[20756] <= 3'b111;
      // memory_array[20757] <= 3'b111;
      // memory_array[20758] <= 3'b111;
      // memory_array[20759] <= 3'b111;
      // memory_array[20760] <= 3'b000;
      // memory_array[20761] <= 3'b000;
      // memory_array[20762] <= 3'b111;
      // memory_array[20763] <= 3'b111;
      // memory_array[20764] <= 3'b111;
      // memory_array[20765] <= 3'b111;
      // memory_array[20766] <= 3'b110;
      // memory_array[20767] <= 3'b000;
      // memory_array[20768] <= 3'b111;
      // memory_array[20769] <= 3'b111;
      // memory_array[20770] <= 3'b111;
      // memory_array[20771] <= 3'b000;
      // memory_array[20772] <= 3'b000;
      // memory_array[20773] <= 3'b111;
      // memory_array[20774] <= 3'b000;
      // memory_array[20775] <= 3'b111;
      // memory_array[20776] <= 3'b111;
      // memory_array[20777] <= 3'b111;
      // memory_array[20778] <= 3'b111;
      // memory_array[20779] <= 3'b110;
      // memory_array[20780] <= 3'b110;
      // memory_array[20781] <= 3'b110;
      // memory_array[20782] <= 3'b110;
      // memory_array[20783] <= 3'b000;
      // memory_array[20784] <= 3'b000;
      // memory_array[20785] <= 3'b110;
      // memory_array[20786] <= 3'b110;
      // memory_array[20787] <= 3'b110;
      // memory_array[20788] <= 3'b000;
      // memory_array[20789] <= 3'b000;
      // memory_array[20790] <= 3'b000;
      // memory_array[20791] <= 3'b101;
      // memory_array[20792] <= 3'b101;
      // memory_array[20793] <= 3'b101;
      // memory_array[20794] <= 3'b000;
      // memory_array[20795] <= 3'b101;
      // memory_array[20796] <= 3'b101;
      // memory_array[20797] <= 3'b110;
      // memory_array[20798] <= 3'b101;
      // memory_array[20799] <= 3'b101;
      // memory_array[20800] <= 3'b101;
      // memory_array[20801] <= 3'b110;
      // memory_array[20802] <= 3'b110;
      // memory_array[20803] <= 3'b000;
      // memory_array[20804] <= 3'b000;
      // memory_array[20805] <= 3'b110;
      // memory_array[20806] <= 3'b110;
      // memory_array[20807] <= 3'b101;
      // memory_array[20808] <= 3'b101;
      // memory_array[20809] <= 3'b000;
      // memory_array[20810] <= 3'b000;
      // memory_array[20811] <= 3'b110;
      // memory_array[20812] <= 3'b110;
      // memory_array[20813] <= 3'b110;
      // memory_array[20814] <= 3'b110;
      // memory_array[20815] <= 3'b110;
      // memory_array[20816] <= 3'b110;
      // memory_array[20817] <= 3'b110;
      // memory_array[20818] <= 3'b111;
      // memory_array[20819] <= 3'b111;
      // memory_array[20820] <= 3'b110;
      // memory_array[20821] <= 3'b000;
      // memory_array[20822] <= 3'b110;
      // memory_array[20823] <= 3'b000;
      // memory_array[20824] <= 3'b111;
      // memory_array[20825] <= 3'b111;
      // memory_array[20826] <= 3'b111;
      // memory_array[20827] <= 3'b111;
      // memory_array[20828] <= 3'b000;
      // memory_array[20829] <= 3'b111;
      // memory_array[20830] <= 3'b111;
      // memory_array[20831] <= 3'b111;
      // memory_array[20832] <= 3'b111;
      // memory_array[20833] <= 3'b000;
      // memory_array[20834] <= 3'b110;
      // memory_array[20835] <= 3'b110;
      // memory_array[20836] <= 3'b110;
      // memory_array[20837] <= 3'b111;
      // memory_array[20838] <= 3'b111;
      // memory_array[20839] <= 3'b111;
      // memory_array[20840] <= 3'b111;
      // memory_array[20841] <= 3'b111;
      // memory_array[20842] <= 3'b111;
      // memory_array[20843] <= 3'b111;
      // memory_array[20844] <= 3'b111;
      // memory_array[20845] <= 3'b000;
      // memory_array[20846] <= 3'b111;
      // memory_array[20847] <= 3'b111;
      // memory_array[20848] <= 3'b111;
      // memory_array[20849] <= 3'b101;
      // memory_array[20850] <= 3'b000;
      // memory_array[20851] <= 3'b111;
      // memory_array[20852] <= 3'b111;
      // memory_array[20853] <= 3'b111;
      // memory_array[20854] <= 3'b111;
      // memory_array[20855] <= 3'b000;
      // memory_array[20856] <= 3'b101;
      // memory_array[20857] <= 3'b111;
      // memory_array[20858] <= 3'b111;
      // memory_array[20859] <= 3'b111;
      // memory_array[20860] <= 3'b111;
      // memory_array[20861] <= 3'b000;
      // memory_array[20862] <= 3'b000;
      // memory_array[20863] <= 3'b000;
      // memory_array[20864] <= 3'b000;
      // memory_array[20865] <= 3'b101;
      // memory_array[20866] <= 3'b101;
      // memory_array[20867] <= 3'b111;
      // memory_array[20868] <= 3'b111;
      // memory_array[20869] <= 3'b111;
      // memory_array[20870] <= 3'b111;
      // memory_array[20871] <= 3'b000;
      // memory_array[20872] <= 3'b101;
      // memory_array[20873] <= 3'b000;
      // memory_array[20874] <= 3'b111;
      // memory_array[20875] <= 3'b111;
      // memory_array[20876] <= 3'b111;
      // memory_array[20877] <= 3'b111;
      // memory_array[20878] <= 3'b000;
      // memory_array[20879] <= 3'b000;
      // memory_array[20880] <= 3'b000;
      // memory_array[20881] <= 3'b000;
      // memory_array[20882] <= 3'b111;
      // memory_array[20883] <= 3'b111;
      // memory_array[20884] <= 3'b111;
      // memory_array[20885] <= 3'b111;
      // memory_array[20886] <= 3'b111;
      // memory_array[20887] <= 3'b111;
      // memory_array[20888] <= 3'b111;
      // memory_array[20889] <= 3'b000;
      // memory_array[20890] <= 3'b000;
      // memory_array[20891] <= 3'b000;
      // memory_array[20892] <= 3'b111;
      // memory_array[20893] <= 3'b111;
      // memory_array[20894] <= 3'b111;
      // memory_array[20895] <= 3'b111;
      // memory_array[20896] <= 3'b000;
      // memory_array[20897] <= 3'b101;
      // memory_array[20898] <= 3'b000;
      // memory_array[20899] <= 3'b000;
      // memory_array[20900] <= 3'b000;
      // memory_array[20901] <= 3'b111;
      // memory_array[20902] <= 3'b111;
      // memory_array[20903] <= 3'b000;
      // memory_array[20904] <= 3'b110;
      // memory_array[20905] <= 3'b110;
      // memory_array[20906] <= 3'b000;
      // memory_array[20907] <= 3'b000;
      // memory_array[20908] <= 3'b111;
      // memory_array[20909] <= 3'b111;
      // memory_array[20910] <= 3'b111;
      // memory_array[20911] <= 3'b111;
      // memory_array[20912] <= 3'b101;
      // memory_array[20913] <= 3'b000;
      // memory_array[20914] <= 3'b101;
      // memory_array[20915] <= 3'b101;
      // memory_array[20916] <= 3'b000;
      // memory_array[20917] <= 3'b000;
      // memory_array[20918] <= 3'b000;
      // memory_array[20919] <= 3'b000;
      // memory_array[20920] <= 3'b000;
      // memory_array[20921] <= 3'b000;
      // memory_array[20922] <= 3'b111;
      // memory_array[20923] <= 3'b111;
      // memory_array[20924] <= 3'b111;
      // memory_array[20925] <= 3'b111;
      // memory_array[20926] <= 3'b111;
      // memory_array[20927] <= 3'b111;
      // memory_array[20928] <= 3'b111;
      // memory_array[20929] <= 3'b111;
      // memory_array[20930] <= 3'b111;
      // memory_array[20931] <= 3'b111;
      // memory_array[20932] <= 3'b111;
      // memory_array[20933] <= 3'b111;
      // memory_array[20934] <= 3'b000;
      // memory_array[20935] <= 3'b111;
      // memory_array[20936] <= 3'b111;
      // memory_array[20937] <= 3'b111;
      // memory_array[20938] <= 3'b111;
      // memory_array[20939] <= 3'b000;
      // memory_array[20940] <= 3'b101;
      // memory_array[20941] <= 3'b111;
      // memory_array[20942] <= 3'b111;
      // memory_array[20943] <= 3'b111;
      // memory_array[20944] <= 3'b111;
      // memory_array[20945] <= 3'b000;
      // memory_array[20946] <= 3'b000;
      // memory_array[20947] <= 3'b000;
      // memory_array[20948] <= 3'b111;
      // memory_array[20949] <= 3'b111;
      // memory_array[20950] <= 3'b111;
      // memory_array[20951] <= 3'b111;
      // memory_array[20952] <= 3'b111;
      // memory_array[20953] <= 3'b000;
      // memory_array[20954] <= 3'b111;
      // memory_array[20955] <= 3'b101;
      // memory_array[20956] <= 3'b111;
      // memory_array[20957] <= 3'b111;
      // memory_array[20958] <= 3'b111;
      // memory_array[20959] <= 3'b111;
      // memory_array[20960] <= 3'b111;
      // memory_array[20961] <= 3'b000;
      // memory_array[20962] <= 3'b111;
      // memory_array[20963] <= 3'b111;
      // memory_array[20964] <= 3'b111;
      // memory_array[20965] <= 3'b111;
      // memory_array[20966] <= 3'b110;
      // memory_array[20967] <= 3'b111;
      // memory_array[20968] <= 3'b111;
      // memory_array[20969] <= 3'b111;
      // memory_array[20970] <= 3'b111;
      // memory_array[20971] <= 3'b110;
      // memory_array[20972] <= 3'b000;
      // memory_array[20973] <= 3'b110;
      // memory_array[20974] <= 3'b000;
      // memory_array[20975] <= 3'b111;
      // memory_array[20976] <= 3'b111;
      // memory_array[20977] <= 3'b111;
      // memory_array[20978] <= 3'b111;
      // memory_array[20979] <= 3'b110;
      // memory_array[20980] <= 3'b110;
      // memory_array[20981] <= 3'b110;
      // memory_array[20982] <= 3'b110;
      // memory_array[20983] <= 3'b111;
      // memory_array[20984] <= 3'b000;
      // memory_array[20985] <= 3'b110;
      // memory_array[20986] <= 3'b110;
      // memory_array[20987] <= 3'b110;
      // memory_array[20988] <= 3'b110;
      // memory_array[20989] <= 3'b000;
      // memory_array[20990] <= 3'b000;
      // memory_array[20991] <= 3'b101;
      // memory_array[20992] <= 3'b110;
      // memory_array[20993] <= 3'b000;
      // memory_array[20994] <= 3'b000;
      // memory_array[20995] <= 3'b110;
      // memory_array[20996] <= 3'b110;
      // memory_array[20997] <= 3'b110;
      // memory_array[20998] <= 3'b000;
      // memory_array[20999] <= 3'b101;
      // memory_array[21000] <= 3'b000;
      // memory_array[21001] <= 3'b000;
      // memory_array[21002] <= 3'b000;
      // memory_array[21003] <= 3'b110;
      // memory_array[21004] <= 3'b110;
      // memory_array[21005] <= 3'b000;
      // memory_array[21006] <= 3'b000;
      // memory_array[21007] <= 3'b000;
      // memory_array[21008] <= 3'b101;
      // memory_array[21009] <= 3'b000;
      // memory_array[21010] <= 3'b000;
      // memory_array[21011] <= 3'b110;
      // memory_array[21012] <= 3'b000;
      // memory_array[21013] <= 3'b110;
      // memory_array[21014] <= 3'b110;
      // memory_array[21015] <= 3'b000;
      // memory_array[21016] <= 3'b111;
      // memory_array[21017] <= 3'b110;
      // memory_array[21018] <= 3'b110;
      // memory_array[21019] <= 3'b110;
      // memory_array[21020] <= 3'b110;
      // memory_array[21021] <= 3'b000;
      // memory_array[21022] <= 3'b111;
      // memory_array[21023] <= 3'b000;
      // memory_array[21024] <= 3'b111;
      // memory_array[21025] <= 3'b111;
      // memory_array[21026] <= 3'b111;
      // memory_array[21027] <= 3'b111;
      // memory_array[21028] <= 3'b111;
      // memory_array[21029] <= 3'b111;
      // memory_array[21030] <= 3'b111;
      // memory_array[21031] <= 3'b111;
      // memory_array[21032] <= 3'b000;
      // memory_array[21033] <= 3'b110;
      // memory_array[21034] <= 3'b110;
      // memory_array[21035] <= 3'b111;
      // memory_array[21036] <= 3'b111;
      // memory_array[21037] <= 3'b111;
      // memory_array[21038] <= 3'b111;
      // memory_array[21039] <= 3'b111;
      // memory_array[21040] <= 3'b111;
      // memory_array[21041] <= 3'b111;
      // memory_array[21042] <= 3'b111;
      // memory_array[21043] <= 3'b111;
      // memory_array[21044] <= 3'b111;
      // memory_array[21045] <= 3'b111;
      // memory_array[21046] <= 3'b111;
      // memory_array[21047] <= 3'b111;
      // memory_array[21048] <= 3'b111;
      // memory_array[21049] <= 3'b101;
      // memory_array[21050] <= 3'b000;
      // memory_array[21051] <= 3'b111;
      // memory_array[21052] <= 3'b111;
      // memory_array[21053] <= 3'b111;
      // memory_array[21054] <= 3'b111;
      // memory_array[21055] <= 3'b000;
      // memory_array[21056] <= 3'b000;
      // memory_array[21057] <= 3'b111;
      // memory_array[21058] <= 3'b111;
      // memory_array[21059] <= 3'b111;
      // memory_array[21060] <= 3'b111;
      // memory_array[21061] <= 3'b000;
      // memory_array[21062] <= 3'b000;
      // memory_array[21063] <= 3'b000;
      // memory_array[21064] <= 3'b000;
      // memory_array[21065] <= 3'b000;
      // memory_array[21066] <= 3'b000;
      // memory_array[21067] <= 3'b111;
      // memory_array[21068] <= 3'b111;
      // memory_array[21069] <= 3'b111;
      // memory_array[21070] <= 3'b111;
      // memory_array[21071] <= 3'b000;
      // memory_array[21072] <= 3'b000;
      // memory_array[21073] <= 3'b000;
      // memory_array[21074] <= 3'b111;
      // memory_array[21075] <= 3'b111;
      // memory_array[21076] <= 3'b111;
      // memory_array[21077] <= 3'b111;
      // memory_array[21078] <= 3'b111;
      // memory_array[21079] <= 3'b000;
      // memory_array[21080] <= 3'b000;
      // memory_array[21081] <= 3'b000;
      // memory_array[21082] <= 3'b111;
      // memory_array[21083] <= 3'b111;
      // memory_array[21084] <= 3'b111;
      // memory_array[21085] <= 3'b111;
      // memory_array[21086] <= 3'b111;
      // memory_array[21087] <= 3'b111;
      // memory_array[21088] <= 3'b111;
      // memory_array[21089] <= 3'b111;
      // memory_array[21090] <= 3'b111;
      // memory_array[21091] <= 3'b111;
      // memory_array[21092] <= 3'b111;
      // memory_array[21093] <= 3'b111;
      // memory_array[21094] <= 3'b000;
      // memory_array[21095] <= 3'b000;
      // memory_array[21096] <= 3'b000;
      // memory_array[21097] <= 3'b000;
      // memory_array[21098] <= 3'b000;
      // memory_array[21099] <= 3'b000;
      // memory_array[21100] <= 3'b000;
      // memory_array[21101] <= 3'b111;
      // memory_array[21102] <= 3'b111;
      // memory_array[21103] <= 3'b000;
      // memory_array[21104] <= 3'b000;
      // memory_array[21105] <= 3'b000;
      // memory_array[21106] <= 3'b000;
      // memory_array[21107] <= 3'b000;
      // memory_array[21108] <= 3'b111;
      // memory_array[21109] <= 3'b111;
      // memory_array[21110] <= 3'b111;
      // memory_array[21111] <= 3'b111;
      // memory_array[21112] <= 3'b000;
      // memory_array[21113] <= 3'b000;
      // memory_array[21114] <= 3'b101;
      // memory_array[21115] <= 3'b000;
      // memory_array[21116] <= 3'b000;
      // memory_array[21117] <= 3'b000;
      // memory_array[21118] <= 3'b000;
      // memory_array[21119] <= 3'b000;
      // memory_array[21120] <= 3'b000;
      // memory_array[21121] <= 3'b000;
      // memory_array[21122] <= 3'b000;
      // memory_array[21123] <= 3'b111;
      // memory_array[21124] <= 3'b111;
      // memory_array[21125] <= 3'b111;
      // memory_array[21126] <= 3'b111;
      // memory_array[21127] <= 3'b111;
      // memory_array[21128] <= 3'b111;
      // memory_array[21129] <= 3'b111;
      // memory_array[21130] <= 3'b111;
      // memory_array[21131] <= 3'b000;
      // memory_array[21132] <= 3'b000;
      // memory_array[21133] <= 3'b000;
      // memory_array[21134] <= 3'b000;
      // memory_array[21135] <= 3'b111;
      // memory_array[21136] <= 3'b111;
      // memory_array[21137] <= 3'b111;
      // memory_array[21138] <= 3'b111;
      // memory_array[21139] <= 3'b101;
      // memory_array[21140] <= 3'b000;
      // memory_array[21141] <= 3'b111;
      // memory_array[21142] <= 3'b111;
      // memory_array[21143] <= 3'b111;
      // memory_array[21144] <= 3'b111;
      // memory_array[21145] <= 3'b000;
      // memory_array[21146] <= 3'b000;
      // memory_array[21147] <= 3'b000;
      // memory_array[21148] <= 3'b000;
      // memory_array[21149] <= 3'b111;
      // memory_array[21150] <= 3'b111;
      // memory_array[21151] <= 3'b111;
      // memory_array[21152] <= 3'b111;
      // memory_array[21153] <= 3'b000;
      // memory_array[21154] <= 3'b111;
      // memory_array[21155] <= 3'b101;
      // memory_array[21156] <= 3'b111;
      // memory_array[21157] <= 3'b111;
      // memory_array[21158] <= 3'b111;
      // memory_array[21159] <= 3'b111;
      // memory_array[21160] <= 3'b111;
      // memory_array[21161] <= 3'b000;
      // memory_array[21162] <= 3'b111;
      // memory_array[21163] <= 3'b111;
      // memory_array[21164] <= 3'b111;
      // memory_array[21165] <= 3'b111;
      // memory_array[21166] <= 3'b110;
      // memory_array[21167] <= 3'b111;
      // memory_array[21168] <= 3'b111;
      // memory_array[21169] <= 3'b111;
      // memory_array[21170] <= 3'b111;
      // memory_array[21171] <= 3'b111;
      // memory_array[21172] <= 3'b000;
      // memory_array[21173] <= 3'b110;
      // memory_array[21174] <= 3'b000;
      // memory_array[21175] <= 3'b111;
      // memory_array[21176] <= 3'b111;
      // memory_array[21177] <= 3'b111;
      // memory_array[21178] <= 3'b111;
      // memory_array[21179] <= 3'b110;
      // memory_array[21180] <= 3'b111;
      // memory_array[21181] <= 3'b111;
      // memory_array[21182] <= 3'b111;
      // memory_array[21183] <= 3'b110;
      // memory_array[21184] <= 3'b110;
      // memory_array[21185] <= 3'b000;
      // memory_array[21186] <= 3'b000;
      // memory_array[21187] <= 3'b000;
      // memory_array[21188] <= 3'b110;
      // memory_array[21189] <= 3'b000;
      // memory_array[21190] <= 3'b000;
      // memory_array[21191] <= 3'b101;
      // memory_array[21192] <= 3'b000;
      // memory_array[21193] <= 3'b110;
      // memory_array[21194] <= 3'b110;
      // memory_array[21195] <= 3'b000;
      // memory_array[21196] <= 3'b000;
      // memory_array[21197] <= 3'b000;
      // memory_array[21198] <= 3'b110;
      // memory_array[21199] <= 3'b110;
      // memory_array[21200] <= 3'b101;
      // memory_array[21201] <= 3'b101;
      // memory_array[21202] <= 3'b101;
      // memory_array[21203] <= 3'b101;
      // memory_array[21204] <= 3'b101;
      // memory_array[21205] <= 3'b101;
      // memory_array[21206] <= 3'b101;
      // memory_array[21207] <= 3'b101;
      // memory_array[21208] <= 3'b101;
      // memory_array[21209] <= 3'b000;
      // memory_array[21210] <= 3'b000;
      // memory_array[21211] <= 3'b110;
      // memory_array[21212] <= 3'b110;
      // memory_array[21213] <= 3'b000;
      // memory_array[21214] <= 3'b000;
      // memory_array[21215] <= 3'b110;
      // memory_array[21216] <= 3'b110;
      // memory_array[21217] <= 3'b110;
      // memory_array[21218] <= 3'b110;
      // memory_array[21219] <= 3'b110;
      // memory_array[21220] <= 3'b110;
      // memory_array[21221] <= 3'b000;
      // memory_array[21222] <= 3'b110;
      // memory_array[21223] <= 3'b000;
      // memory_array[21224] <= 3'b111;
      // memory_array[21225] <= 3'b111;
      // memory_array[21226] <= 3'b111;
      // memory_array[21227] <= 3'b111;
      // memory_array[21228] <= 3'b111;
      // memory_array[21229] <= 3'b111;
      // memory_array[21230] <= 3'b111;
      // memory_array[21231] <= 3'b000;
      // memory_array[21232] <= 3'b000;
      // memory_array[21233] <= 3'b110;
      // memory_array[21234] <= 3'b111;
      // memory_array[21235] <= 3'b110;
      // memory_array[21236] <= 3'b110;
      // memory_array[21237] <= 3'b111;
      // memory_array[21238] <= 3'b111;
      // memory_array[21239] <= 3'b111;
      // memory_array[21240] <= 3'b111;
      // memory_array[21241] <= 3'b111;
      // memory_array[21242] <= 3'b111;
      // memory_array[21243] <= 3'b111;
      // memory_array[21244] <= 3'b111;
      // memory_array[21245] <= 3'b111;
      // memory_array[21246] <= 3'b111;
      // memory_array[21247] <= 3'b111;
      // memory_array[21248] <= 3'b111;
      // memory_array[21249] <= 3'b101;
      // memory_array[21250] <= 3'b000;
      // memory_array[21251] <= 3'b111;
      // memory_array[21252] <= 3'b111;
      // memory_array[21253] <= 3'b111;
      // memory_array[21254] <= 3'b111;
      // memory_array[21255] <= 3'b000;
      // memory_array[21256] <= 3'b101;
      // memory_array[21257] <= 3'b111;
      // memory_array[21258] <= 3'b111;
      // memory_array[21259] <= 3'b111;
      // memory_array[21260] <= 3'b111;
      // memory_array[21261] <= 3'b000;
      // memory_array[21262] <= 3'b000;
      // memory_array[21263] <= 3'b000;
      // memory_array[21264] <= 3'b000;
      // memory_array[21265] <= 3'b101;
      // memory_array[21266] <= 3'b101;
      // memory_array[21267] <= 3'b111;
      // memory_array[21268] <= 3'b111;
      // memory_array[21269] <= 3'b111;
      // memory_array[21270] <= 3'b111;
      // memory_array[21271] <= 3'b000;
      // memory_array[21272] <= 3'b000;
      // memory_array[21273] <= 3'b000;
      // memory_array[21274] <= 3'b111;
      // memory_array[21275] <= 3'b111;
      // memory_array[21276] <= 3'b111;
      // memory_array[21277] <= 3'b111;
      // memory_array[21278] <= 3'b111;
      // memory_array[21279] <= 3'b000;
      // memory_array[21280] <= 3'b000;
      // memory_array[21281] <= 3'b111;
      // memory_array[21282] <= 3'b111;
      // memory_array[21283] <= 3'b111;
      // memory_array[21284] <= 3'b111;
      // memory_array[21285] <= 3'b111;
      // memory_array[21286] <= 3'b111;
      // memory_array[21287] <= 3'b111;
      // memory_array[21288] <= 3'b111;
      // memory_array[21289] <= 3'b111;
      // memory_array[21290] <= 3'b111;
      // memory_array[21291] <= 3'b111;
      // memory_array[21292] <= 3'b000;
      // memory_array[21293] <= 3'b000;
      // memory_array[21294] <= 3'b000;
      // memory_array[21295] <= 3'b000;
      // memory_array[21296] <= 3'b111;
      // memory_array[21297] <= 3'b000;
      // memory_array[21298] <= 3'b000;
      // memory_array[21299] <= 3'b000;
      // memory_array[21300] <= 3'b000;
      // memory_array[21301] <= 3'b111;
      // memory_array[21302] <= 3'b111;
      // memory_array[21303] <= 3'b000;
      // memory_array[21304] <= 3'b000;
      // memory_array[21305] <= 3'b000;
      // memory_array[21306] <= 3'b101;
      // memory_array[21307] <= 3'b000;
      // memory_array[21308] <= 3'b111;
      // memory_array[21309] <= 3'b111;
      // memory_array[21310] <= 3'b111;
      // memory_array[21311] <= 3'b111;
      // memory_array[21312] <= 3'b000;
      // memory_array[21313] <= 3'b101;
      // memory_array[21314] <= 3'b000;
      // memory_array[21315] <= 3'b101;
      // memory_array[21316] <= 3'b000;
      // memory_array[21317] <= 3'b101;
      // memory_array[21318] <= 3'b000;
      // memory_array[21319] <= 3'b000;
      // memory_array[21320] <= 3'b000;
      // memory_array[21321] <= 3'b000;
      // memory_array[21322] <= 3'b000;
      // memory_array[21323] <= 3'b111;
      // memory_array[21324] <= 3'b111;
      // memory_array[21325] <= 3'b111;
      // memory_array[21326] <= 3'b111;
      // memory_array[21327] <= 3'b111;
      // memory_array[21328] <= 3'b111;
      // memory_array[21329] <= 3'b000;
      // memory_array[21330] <= 3'b000;
      // memory_array[21331] <= 3'b110;
      // memory_array[21332] <= 3'b101;
      // memory_array[21333] <= 3'b000;
      // memory_array[21334] <= 3'b000;
      // memory_array[21335] <= 3'b111;
      // memory_array[21336] <= 3'b111;
      // memory_array[21337] <= 3'b111;
      // memory_array[21338] <= 3'b111;
      // memory_array[21339] <= 3'b000;
      // memory_array[21340] <= 3'b000;
      // memory_array[21341] <= 3'b111;
      // memory_array[21342] <= 3'b111;
      // memory_array[21343] <= 3'b111;
      // memory_array[21344] <= 3'b111;
      // memory_array[21345] <= 3'b111;
      // memory_array[21346] <= 3'b000;
      // memory_array[21347] <= 3'b000;
      // memory_array[21348] <= 3'b000;
      // memory_array[21349] <= 3'b111;
      // memory_array[21350] <= 3'b111;
      // memory_array[21351] <= 3'b111;
      // memory_array[21352] <= 3'b111;
      // memory_array[21353] <= 3'b000;
      // memory_array[21354] <= 3'b111;
      // memory_array[21355] <= 3'b101;
      // memory_array[21356] <= 3'b111;
      // memory_array[21357] <= 3'b111;
      // memory_array[21358] <= 3'b111;
      // memory_array[21359] <= 3'b111;
      // memory_array[21360] <= 3'b111;
      // memory_array[21361] <= 3'b000;
      // memory_array[21362] <= 3'b111;
      // memory_array[21363] <= 3'b111;
      // memory_array[21364] <= 3'b111;
      // memory_array[21365] <= 3'b111;
      // memory_array[21366] <= 3'b000;
      // memory_array[21367] <= 3'b111;
      // memory_array[21368] <= 3'b111;
      // memory_array[21369] <= 3'b111;
      // memory_array[21370] <= 3'b111;
      // memory_array[21371] <= 3'b110;
      // memory_array[21372] <= 3'b000;
      // memory_array[21373] <= 3'b111;
      // memory_array[21374] <= 3'b000;
      // memory_array[21375] <= 3'b111;
      // memory_array[21376] <= 3'b111;
      // memory_array[21377] <= 3'b111;
      // memory_array[21378] <= 3'b111;
      // memory_array[21379] <= 3'b111;
      // memory_array[21380] <= 3'b110;
      // memory_array[21381] <= 3'b110;
      // memory_array[21382] <= 3'b110;
      // memory_array[21383] <= 3'b110;
      // memory_array[21384] <= 3'b110;
      // memory_array[21385] <= 3'b110;
      // memory_array[21386] <= 3'b110;
      // memory_array[21387] <= 3'b110;
      // memory_array[21388] <= 3'b000;
      // memory_array[21389] <= 3'b000;
      // memory_array[21390] <= 3'b000;
      // memory_array[21391] <= 3'b101;
      // memory_array[21392] <= 3'b101;
      // memory_array[21393] <= 3'b101;
      // memory_array[21394] <= 3'b101;
      // memory_array[21395] <= 3'b101;
      // memory_array[21396] <= 3'b101;
      // memory_array[21397] <= 3'b101;
      // memory_array[21398] <= 3'b101;
      // memory_array[21399] <= 3'b101;
      // memory_array[21400] <= 3'b101;
      // memory_array[21401] <= 3'b101;
      // memory_array[21402] <= 3'b101;
      // memory_array[21403] <= 3'b101;
      // memory_array[21404] <= 3'b101;
      // memory_array[21405] <= 3'b101;
      // memory_array[21406] <= 3'b101;
      // memory_array[21407] <= 3'b101;
      // memory_array[21408] <= 3'b101;
      // memory_array[21409] <= 3'b000;
      // memory_array[21410] <= 3'b000;
      // memory_array[21411] <= 3'b110;
      // memory_array[21412] <= 3'b110;
      // memory_array[21413] <= 3'b000;
      // memory_array[21414] <= 3'b000;
      // memory_array[21415] <= 3'b110;
      // memory_array[21416] <= 3'b110;
      // memory_array[21417] <= 3'b110;
      // memory_array[21418] <= 3'b110;
      // memory_array[21419] <= 3'b110;
      // memory_array[21420] <= 3'b110;
      // memory_array[21421] <= 3'b000;
      // memory_array[21422] <= 3'b110;
      // memory_array[21423] <= 3'b000;
      // memory_array[21424] <= 3'b111;
      // memory_array[21425] <= 3'b111;
      // memory_array[21426] <= 3'b111;
      // memory_array[21427] <= 3'b000;
      // memory_array[21428] <= 3'b000;
      // memory_array[21429] <= 3'b000;
      // memory_array[21430] <= 3'b110;
      // memory_array[21431] <= 3'b110;
      // memory_array[21432] <= 3'b000;
      // memory_array[21433] <= 3'b110;
      // memory_array[21434] <= 3'b111;
      // memory_array[21435] <= 3'b110;
      // memory_array[21436] <= 3'b110;
      // memory_array[21437] <= 3'b111;
      // memory_array[21438] <= 3'b111;
      // memory_array[21439] <= 3'b111;
      // memory_array[21440] <= 3'b111;
      // memory_array[21441] <= 3'b000;
      // memory_array[21442] <= 3'b111;
      // memory_array[21443] <= 3'b111;
      // memory_array[21444] <= 3'b111;
      // memory_array[21445] <= 3'b111;
      // memory_array[21446] <= 3'b000;
      // memory_array[21447] <= 3'b111;
      // memory_array[21448] <= 3'b111;
      // memory_array[21449] <= 3'b101;
      // memory_array[21450] <= 3'b000;
      // memory_array[21451] <= 3'b111;
      // memory_array[21452] <= 3'b111;
      // memory_array[21453] <= 3'b111;
      // memory_array[21454] <= 3'b111;
      // memory_array[21455] <= 3'b000;
      // memory_array[21456] <= 3'b101;
      // memory_array[21457] <= 3'b111;
      // memory_array[21458] <= 3'b111;
      // memory_array[21459] <= 3'b111;
      // memory_array[21460] <= 3'b111;
      // memory_array[21461] <= 3'b000;
      // memory_array[21462] <= 3'b101;
      // memory_array[21463] <= 3'b000;
      // memory_array[21464] <= 3'b000;
      // memory_array[21465] <= 3'b000;
      // memory_array[21466] <= 3'b101;
      // memory_array[21467] <= 3'b111;
      // memory_array[21468] <= 3'b111;
      // memory_array[21469] <= 3'b111;
      // memory_array[21470] <= 3'b111;
      // memory_array[21471] <= 3'b000;
      // memory_array[21472] <= 3'b000;
      // memory_array[21473] <= 3'b000;
      // memory_array[21474] <= 3'b000;
      // memory_array[21475] <= 3'b000;
      // memory_array[21476] <= 3'b111;
      // memory_array[21477] <= 3'b111;
      // memory_array[21478] <= 3'b111;
      // memory_array[21479] <= 3'b111;
      // memory_array[21480] <= 3'b111;
      // memory_array[21481] <= 3'b111;
      // memory_array[21482] <= 3'b111;
      // memory_array[21483] <= 3'b111;
      // memory_array[21484] <= 3'b000;
      // memory_array[21485] <= 3'b000;
      // memory_array[21486] <= 3'b111;
      // memory_array[21487] <= 3'b111;
      // memory_array[21488] <= 3'b000;
      // memory_array[21489] <= 3'b000;
      // memory_array[21490] <= 3'b000;
      // memory_array[21491] <= 3'b000;
      // memory_array[21492] <= 3'b111;
      // memory_array[21493] <= 3'b111;
      // memory_array[21494] <= 3'b111;
      // memory_array[21495] <= 3'b111;
      // memory_array[21496] <= 3'b000;
      // memory_array[21497] <= 3'b000;
      // memory_array[21498] <= 3'b000;
      // memory_array[21499] <= 3'b111;
      // memory_array[21500] <= 3'b111;
      // memory_array[21501] <= 3'b111;
      // memory_array[21502] <= 3'b000;
      // memory_array[21503] <= 3'b000;
      // memory_array[21504] <= 3'b000;
      // memory_array[21505] <= 3'b000;
      // memory_array[21506] <= 3'b000;
      // memory_array[21507] <= 3'b000;
      // memory_array[21508] <= 3'b111;
      // memory_array[21509] <= 3'b111;
      // memory_array[21510] <= 3'b111;
      // memory_array[21511] <= 3'b111;
      // memory_array[21512] <= 3'b111;
      // memory_array[21513] <= 3'b000;
      // memory_array[21514] <= 3'b000;
      // memory_array[21515] <= 3'b000;
      // memory_array[21516] <= 3'b000;
      // memory_array[21517] <= 3'b101;
      // memory_array[21518] <= 3'b000;
      // memory_array[21519] <= 3'b000;
      // memory_array[21520] <= 3'b000;
      // memory_array[21521] <= 3'b000;
      // memory_array[21522] <= 3'b101;
      // memory_array[21523] <= 3'b000;
      // memory_array[21524] <= 3'b111;
      // memory_array[21525] <= 3'b111;
      // memory_array[21526] <= 3'b111;
      // memory_array[21527] <= 3'b000;
      // memory_array[21528] <= 3'b000;
      // memory_array[21529] <= 3'b000;
      // memory_array[21530] <= 3'b000;
      // memory_array[21531] <= 3'b101;
      // memory_array[21532] <= 3'b101;
      // memory_array[21533] <= 3'b000;
      // memory_array[21534] <= 3'b000;
      // memory_array[21535] <= 3'b111;
      // memory_array[21536] <= 3'b111;
      // memory_array[21537] <= 3'b111;
      // memory_array[21538] <= 3'b111;
      // memory_array[21539] <= 3'b000;
      // memory_array[21540] <= 3'b000;
      // memory_array[21541] <= 3'b000;
      // memory_array[21542] <= 3'b111;
      // memory_array[21543] <= 3'b111;
      // memory_array[21544] <= 3'b111;
      // memory_array[21545] <= 3'b111;
      // memory_array[21546] <= 3'b000;
      // memory_array[21547] <= 3'b000;
      // memory_array[21548] <= 3'b111;
      // memory_array[21549] <= 3'b111;
      // memory_array[21550] <= 3'b111;
      // memory_array[21551] <= 3'b111;
      // memory_array[21552] <= 3'b000;
      // memory_array[21553] <= 3'b111;
      // memory_array[21554] <= 3'b111;
      // memory_array[21555] <= 3'b101;
      // memory_array[21556] <= 3'b111;
      // memory_array[21557] <= 3'b111;
      // memory_array[21558] <= 3'b111;
      // memory_array[21559] <= 3'b111;
      // memory_array[21560] <= 3'b111;
      // memory_array[21561] <= 3'b000;
      // memory_array[21562] <= 3'b111;
      // memory_array[21563] <= 3'b111;
      // memory_array[21564] <= 3'b111;
      // memory_array[21565] <= 3'b111;
      // memory_array[21566] <= 3'b000;
      // memory_array[21567] <= 3'b111;
      // memory_array[21568] <= 3'b111;
      // memory_array[21569] <= 3'b111;
      // memory_array[21570] <= 3'b111;
      // memory_array[21571] <= 3'b110;
      // memory_array[21572] <= 3'b000;
      // memory_array[21573] <= 3'b111;
      // memory_array[21574] <= 3'b000;
      // memory_array[21575] <= 3'b111;
      // memory_array[21576] <= 3'b111;
      // memory_array[21577] <= 3'b111;
      // memory_array[21578] <= 3'b111;
      // memory_array[21579] <= 3'b111;
      // memory_array[21580] <= 3'b110;
      // memory_array[21581] <= 3'b110;
      // memory_array[21582] <= 3'b110;
      // memory_array[21583] <= 3'b110;
      // memory_array[21584] <= 3'b110;
      // memory_array[21585] <= 3'b110;
      // memory_array[21586] <= 3'b110;
      // memory_array[21587] <= 3'b110;
      // memory_array[21588] <= 3'b000;
      // memory_array[21589] <= 3'b000;
      // memory_array[21590] <= 3'b000;
      // memory_array[21591] <= 3'b101;
      // memory_array[21592] <= 3'b101;
      // memory_array[21593] <= 3'b101;
      // memory_array[21594] <= 3'b101;
      // memory_array[21595] <= 3'b101;
      // memory_array[21596] <= 3'b101;
      // memory_array[21597] <= 3'b101;
      // memory_array[21598] <= 3'b101;
      // memory_array[21599] <= 3'b101;
      // memory_array[21600] <= 3'b000;
      // memory_array[21601] <= 3'b000;
      // memory_array[21602] <= 3'b000;
      // memory_array[21603] <= 3'b110;
      // memory_array[21604] <= 3'b110;
      // memory_array[21605] <= 3'b000;
      // memory_array[21606] <= 3'b000;
      // memory_array[21607] <= 3'b000;
      // memory_array[21608] <= 3'b101;
      // memory_array[21609] <= 3'b000;
      // memory_array[21610] <= 3'b000;
      // memory_array[21611] <= 3'b110;
      // memory_array[21612] <= 3'b000;
      // memory_array[21613] <= 3'b110;
      // memory_array[21614] <= 3'b110;
      // memory_array[21615] <= 3'b000;
      // memory_array[21616] <= 3'b111;
      // memory_array[21617] <= 3'b110;
      // memory_array[21618] <= 3'b110;
      // memory_array[21619] <= 3'b110;
      // memory_array[21620] <= 3'b110;
      // memory_array[21621] <= 3'b000;
      // memory_array[21622] <= 3'b111;
      // memory_array[21623] <= 3'b000;
      // memory_array[21624] <= 3'b111;
      // memory_array[21625] <= 3'b111;
      // memory_array[21626] <= 3'b111;
      // memory_array[21627] <= 3'b000;
      // memory_array[21628] <= 3'b110;
      // memory_array[21629] <= 3'b110;
      // memory_array[21630] <= 3'b110;
      // memory_array[21631] <= 3'b110;
      // memory_array[21632] <= 3'b000;
      // memory_array[21633] <= 3'b110;
      // memory_array[21634] <= 3'b110;
      // memory_array[21635] <= 3'b111;
      // memory_array[21636] <= 3'b111;
      // memory_array[21637] <= 3'b111;
      // memory_array[21638] <= 3'b111;
      // memory_array[21639] <= 3'b111;
      // memory_array[21640] <= 3'b111;
      // memory_array[21641] <= 3'b000;
      // memory_array[21642] <= 3'b111;
      // memory_array[21643] <= 3'b111;
      // memory_array[21644] <= 3'b111;
      // memory_array[21645] <= 3'b111;
      // memory_array[21646] <= 3'b111;
      // memory_array[21647] <= 3'b111;
      // memory_array[21648] <= 3'b111;
      // memory_array[21649] <= 3'b101;
      // memory_array[21650] <= 3'b000;
      // memory_array[21651] <= 3'b111;
      // memory_array[21652] <= 3'b111;
      // memory_array[21653] <= 3'b111;
      // memory_array[21654] <= 3'b111;
      // memory_array[21655] <= 3'b000;
      // memory_array[21656] <= 3'b000;
      // memory_array[21657] <= 3'b111;
      // memory_array[21658] <= 3'b111;
      // memory_array[21659] <= 3'b111;
      // memory_array[21660] <= 3'b111;
      // memory_array[21661] <= 3'b000;
      // memory_array[21662] <= 3'b000;
      // memory_array[21663] <= 3'b101;
      // memory_array[21664] <= 3'b101;
      // memory_array[21665] <= 3'b000;
      // memory_array[21666] <= 3'b000;
      // memory_array[21667] <= 3'b111;
      // memory_array[21668] <= 3'b111;
      // memory_array[21669] <= 3'b111;
      // memory_array[21670] <= 3'b111;
      // memory_array[21671] <= 3'b111;
      // memory_array[21672] <= 3'b000;
      // memory_array[21673] <= 3'b000;
      // memory_array[21674] <= 3'b000;
      // memory_array[21675] <= 3'b000;
      // memory_array[21676] <= 3'b000;
      // memory_array[21677] <= 3'b111;
      // memory_array[21678] <= 3'b111;
      // memory_array[21679] <= 3'b111;
      // memory_array[21680] <= 3'b111;
      // memory_array[21681] <= 3'b111;
      // memory_array[21682] <= 3'b000;
      // memory_array[21683] <= 3'b000;
      // memory_array[21684] <= 3'b101;
      // memory_array[21685] <= 3'b000;
      // memory_array[21686] <= 3'b000;
      // memory_array[21687] <= 3'b000;
      // memory_array[21688] <= 3'b000;
      // memory_array[21689] <= 3'b000;
      // memory_array[21690] <= 3'b000;
      // memory_array[21691] <= 3'b111;
      // memory_array[21692] <= 3'b111;
      // memory_array[21693] <= 3'b111;
      // memory_array[21694] <= 3'b111;
      // memory_array[21695] <= 3'b111;
      // memory_array[21696] <= 3'b111;
      // memory_array[21697] <= 3'b111;
      // memory_array[21698] <= 3'b111;
      // memory_array[21699] <= 3'b111;
      // memory_array[21700] <= 3'b111;
      // memory_array[21701] <= 3'b111;
      // memory_array[21702] <= 3'b000;
      // memory_array[21703] <= 3'b000;
      // memory_array[21704] <= 3'b000;
      // memory_array[21705] <= 3'b000;
      // memory_array[21706] <= 3'b000;
      // memory_array[21707] <= 3'b111;
      // memory_array[21708] <= 3'b111;
      // memory_array[21709] <= 3'b111;
      // memory_array[21710] <= 3'b111;
      // memory_array[21711] <= 3'b000;
      // memory_array[21712] <= 3'b000;
      // memory_array[21713] <= 3'b000;
      // memory_array[21714] <= 3'b101;
      // memory_array[21715] <= 3'b000;
      // memory_array[21716] <= 3'b000;
      // memory_array[21717] <= 3'b000;
      // memory_array[21718] <= 3'b000;
      // memory_array[21719] <= 3'b101;
      // memory_array[21720] <= 3'b000;
      // memory_array[21721] <= 3'b000;
      // memory_array[21722] <= 3'b000;
      // memory_array[21723] <= 3'b101;
      // memory_array[21724] <= 3'b111;
      // memory_array[21725] <= 3'b111;
      // memory_array[21726] <= 3'b000;
      // memory_array[21727] <= 3'b000;
      // memory_array[21728] <= 3'b101;
      // memory_array[21729] <= 3'b101;
      // memory_array[21730] <= 3'b000;
      // memory_array[21731] <= 3'b000;
      // memory_array[21732] <= 3'b000;
      // memory_array[21733] <= 3'b000;
      // memory_array[21734] <= 3'b000;
      // memory_array[21735] <= 3'b111;
      // memory_array[21736] <= 3'b111;
      // memory_array[21737] <= 3'b111;
      // memory_array[21738] <= 3'b111;
      // memory_array[21739] <= 3'b000;
      // memory_array[21740] <= 3'b000;
      // memory_array[21741] <= 3'b000;
      // memory_array[21742] <= 3'b111;
      // memory_array[21743] <= 3'b111;
      // memory_array[21744] <= 3'b111;
      // memory_array[21745] <= 3'b111;
      // memory_array[21746] <= 3'b000;
      // memory_array[21747] <= 3'b000;
      // memory_array[21748] <= 3'b111;
      // memory_array[21749] <= 3'b111;
      // memory_array[21750] <= 3'b111;
      // memory_array[21751] <= 3'b111;
      // memory_array[21752] <= 3'b111;
      // memory_array[21753] <= 3'b111;
      // memory_array[21754] <= 3'b111;
      // memory_array[21755] <= 3'b101;
      // memory_array[21756] <= 3'b111;
      // memory_array[21757] <= 3'b111;
      // memory_array[21758] <= 3'b111;
      // memory_array[21759] <= 3'b111;
      // memory_array[21760] <= 3'b111;
      // memory_array[21761] <= 3'b000;
      // memory_array[21762] <= 3'b111;
      // memory_array[21763] <= 3'b111;
      // memory_array[21764] <= 3'b111;
      // memory_array[21765] <= 3'b111;
      // memory_array[21766] <= 3'b111;
      // memory_array[21767] <= 3'b111;
      // memory_array[21768] <= 3'b111;
      // memory_array[21769] <= 3'b111;
      // memory_array[21770] <= 3'b111;
      // memory_array[21771] <= 3'b111;
      // memory_array[21772] <= 3'b000;
      // memory_array[21773] <= 3'b110;
      // memory_array[21774] <= 3'b000;
      // memory_array[21775] <= 3'b111;
      // memory_array[21776] <= 3'b111;
      // memory_array[21777] <= 3'b111;
      // memory_array[21778] <= 3'b111;
      // memory_array[21779] <= 3'b110;
      // memory_array[21780] <= 3'b111;
      // memory_array[21781] <= 3'b111;
      // memory_array[21782] <= 3'b111;
      // memory_array[21783] <= 3'b110;
      // memory_array[21784] <= 3'b110;
      // memory_array[21785] <= 3'b000;
      // memory_array[21786] <= 3'b000;
      // memory_array[21787] <= 3'b000;
      // memory_array[21788] <= 3'b110;
      // memory_array[21789] <= 3'b000;
      // memory_array[21790] <= 3'b000;
      // memory_array[21791] <= 3'b101;
      // memory_array[21792] <= 3'b000;
      // memory_array[21793] <= 3'b110;
      // memory_array[21794] <= 3'b110;
      // memory_array[21795] <= 3'b000;
      // memory_array[21796] <= 3'b000;
      // memory_array[21797] <= 3'b000;
      // memory_array[21798] <= 3'b110;
      // memory_array[21799] <= 3'b110;
      // memory_array[21800] <= 3'b101;
      // memory_array[21801] <= 3'b000;
      // memory_array[21802] <= 3'b000;
      // memory_array[21803] <= 3'b110;
      // memory_array[21804] <= 3'b110;
      // memory_array[21805] <= 3'b000;
      // memory_array[21806] <= 3'b000;
      // memory_array[21807] <= 3'b101;
      // memory_array[21808] <= 3'b101;
      // memory_array[21809] <= 3'b000;
      // memory_array[21810] <= 3'b000;
      // memory_array[21811] <= 3'b000;
      // memory_array[21812] <= 3'b000;
      // memory_array[21813] <= 3'b000;
      // memory_array[21814] <= 3'b000;
      // memory_array[21815] <= 3'b000;
      // memory_array[21816] <= 3'b000;
      // memory_array[21817] <= 3'b000;
      // memory_array[21818] <= 3'b000;
      // memory_array[21819] <= 3'b000;
      // memory_array[21820] <= 3'b000;
      // memory_array[21821] <= 3'b000;
      // memory_array[21822] <= 3'b000;
      // memory_array[21823] <= 3'b000;
      // memory_array[21824] <= 3'b111;
      // memory_array[21825] <= 3'b111;
      // memory_array[21826] <= 3'b111;
      // memory_array[21827] <= 3'b000;
      // memory_array[21828] <= 3'b000;
      // memory_array[21829] <= 3'b000;
      // memory_array[21830] <= 3'b000;
      // memory_array[21831] <= 3'b000;
      // memory_array[21832] <= 3'b000;
      // memory_array[21833] <= 3'b000;
      // memory_array[21834] <= 3'b000;
      // memory_array[21835] <= 3'b000;
      // memory_array[21836] <= 3'b000;
      // memory_array[21837] <= 3'b111;
      // memory_array[21838] <= 3'b111;
      // memory_array[21839] <= 3'b111;
      // memory_array[21840] <= 3'b111;
      // memory_array[21841] <= 3'b000;
      // memory_array[21842] <= 3'b000;
      // memory_array[21843] <= 3'b111;
      // memory_array[21844] <= 3'b111;
      // memory_array[21845] <= 3'b111;
      // memory_array[21846] <= 3'b111;
      // memory_array[21847] <= 3'b000;
      // memory_array[21848] <= 3'b111;
      // memory_array[21849] <= 3'b101;
      // memory_array[21850] <= 3'b000;
      // memory_array[21851] <= 3'b111;
      // memory_array[21852] <= 3'b111;
      // memory_array[21853] <= 3'b111;
      // memory_array[21854] <= 3'b111;
      // memory_array[21855] <= 3'b000;
      // memory_array[21856] <= 3'b000;
      // memory_array[21857] <= 3'b111;
      // memory_array[21858] <= 3'b111;
      // memory_array[21859] <= 3'b111;
      // memory_array[21860] <= 3'b111;
      // memory_array[21861] <= 3'b000;
      // memory_array[21862] <= 3'b000;
      // memory_array[21863] <= 3'b000;
      // memory_array[21864] <= 3'b000;
      // memory_array[21865] <= 3'b000;
      // memory_array[21866] <= 3'b000;
      // memory_array[21867] <= 3'b111;
      // memory_array[21868] <= 3'b111;
      // memory_array[21869] <= 3'b111;
      // memory_array[21870] <= 3'b111;
      // memory_array[21871] <= 3'b111;
      // memory_array[21872] <= 3'b000;
      // memory_array[21873] <= 3'b000;
      // memory_array[21874] <= 3'b101;
      // memory_array[21875] <= 3'b000;
      // memory_array[21876] <= 3'b000;
      // memory_array[21877] <= 3'b000;
      // memory_array[21878] <= 3'b101;
      // memory_array[21879] <= 3'b101;
      // memory_array[21880] <= 3'b000;
      // memory_array[21881] <= 3'b101;
      // memory_array[21882] <= 3'b000;
      // memory_array[21883] <= 3'b000;
      // memory_array[21884] <= 3'b101;
      // memory_array[21885] <= 3'b000;
      // memory_array[21886] <= 3'b000;
      // memory_array[21887] <= 3'b000;
      // memory_array[21888] <= 3'b000;
      // memory_array[21889] <= 3'b000;
      // memory_array[21890] <= 3'b000;
      // memory_array[21891] <= 3'b111;
      // memory_array[21892] <= 3'b111;
      // memory_array[21893] <= 3'b111;
      // memory_array[21894] <= 3'b111;
      // memory_array[21895] <= 3'b111;
      // memory_array[21896] <= 3'b111;
      // memory_array[21897] <= 3'b111;
      // memory_array[21898] <= 3'b111;
      // memory_array[21899] <= 3'b000;
      // memory_array[21900] <= 3'b000;
      // memory_array[21901] <= 3'b000;
      // memory_array[21902] <= 3'b000;
      // memory_array[21903] <= 3'b000;
      // memory_array[21904] <= 3'b000;
      // memory_array[21905] <= 3'b000;
      // memory_array[21906] <= 3'b000;
      // memory_array[21907] <= 3'b111;
      // memory_array[21908] <= 3'b000;
      // memory_array[21909] <= 3'b000;
      // memory_array[21910] <= 3'b000;
      // memory_array[21911] <= 3'b000;
      // memory_array[21912] <= 3'b000;
      // memory_array[21913] <= 3'b101;
      // memory_array[21914] <= 3'b101;
      // memory_array[21915] <= 3'b000;
      // memory_array[21916] <= 3'b000;
      // memory_array[21917] <= 3'b000;
      // memory_array[21918] <= 3'b000;
      // memory_array[21919] <= 3'b000;
      // memory_array[21920] <= 3'b000;
      // memory_array[21921] <= 3'b000;
      // memory_array[21922] <= 3'b000;
      // memory_array[21923] <= 3'b101;
      // memory_array[21924] <= 3'b000;
      // memory_array[21925] <= 3'b000;
      // memory_array[21926] <= 3'b000;
      // memory_array[21927] <= 3'b000;
      // memory_array[21928] <= 3'b101;
      // memory_array[21929] <= 3'b101;
      // memory_array[21930] <= 3'b000;
      // memory_array[21931] <= 3'b000;
      // memory_array[21932] <= 3'b000;
      // memory_array[21933] <= 3'b000;
      // memory_array[21934] <= 3'b111;
      // memory_array[21935] <= 3'b111;
      // memory_array[21936] <= 3'b111;
      // memory_array[21937] <= 3'b111;
      // memory_array[21938] <= 3'b111;
      // memory_array[21939] <= 3'b000;
      // memory_array[21940] <= 3'b000;
      // memory_array[21941] <= 3'b000;
      // memory_array[21942] <= 3'b111;
      // memory_array[21943] <= 3'b111;
      // memory_array[21944] <= 3'b111;
      // memory_array[21945] <= 3'b111;
      // memory_array[21946] <= 3'b111;
      // memory_array[21947] <= 3'b000;
      // memory_array[21948] <= 3'b111;
      // memory_array[21949] <= 3'b111;
      // memory_array[21950] <= 3'b111;
      // memory_array[21951] <= 3'b111;
      // memory_array[21952] <= 3'b111;
      // memory_array[21953] <= 3'b111;
      // memory_array[21954] <= 3'b111;
      // memory_array[21955] <= 3'b101;
      // memory_array[21956] <= 3'b111;
      // memory_array[21957] <= 3'b111;
      // memory_array[21958] <= 3'b111;
      // memory_array[21959] <= 3'b111;
      // memory_array[21960] <= 3'b000;
      // memory_array[21961] <= 3'b000;
      // memory_array[21962] <= 3'b111;
      // memory_array[21963] <= 3'b111;
      // memory_array[21964] <= 3'b111;
      // memory_array[21965] <= 3'b111;
      // memory_array[21966] <= 3'b111;
      // memory_array[21967] <= 3'b111;
      // memory_array[21968] <= 3'b111;
      // memory_array[21969] <= 3'b111;
      // memory_array[21970] <= 3'b111;
      // memory_array[21971] <= 3'b000;
      // memory_array[21972] <= 3'b000;
      // memory_array[21973] <= 3'b000;
      // memory_array[21974] <= 3'b000;
      // memory_array[21975] <= 3'b111;
      // memory_array[21976] <= 3'b111;
      // memory_array[21977] <= 3'b111;
      // memory_array[21978] <= 3'b111;
      // memory_array[21979] <= 3'b000;
      // memory_array[21980] <= 3'b000;
      // memory_array[21981] <= 3'b000;
      // memory_array[21982] <= 3'b000;
      // memory_array[21983] <= 3'b000;
      // memory_array[21984] <= 3'b000;
      // memory_array[21985] <= 3'b000;
      // memory_array[21986] <= 3'b000;
      // memory_array[21987] <= 3'b000;
      // memory_array[21988] <= 3'b000;
      // memory_array[21989] <= 3'b000;
      // memory_array[21990] <= 3'b000;
      // memory_array[21991] <= 3'b101;
      // memory_array[21992] <= 3'b101;
      // memory_array[21993] <= 3'b110;
      // memory_array[21994] <= 3'b110;
      // memory_array[21995] <= 3'b000;
      // memory_array[21996] <= 3'b000;
      // memory_array[21997] <= 3'b000;
      // memory_array[21998] <= 3'b110;
      // memory_array[21999] <= 3'b101;
      // memory_array[22000] <= 3'b101;
      // memory_array[22001] <= 3'b000;
      // memory_array[22002] <= 3'b000;
      // memory_array[22003] <= 3'b110;
      // memory_array[22004] <= 3'b110;
      // memory_array[22005] <= 3'b000;
      // memory_array[22006] <= 3'b000;
      // memory_array[22007] <= 3'b101;
      // memory_array[22008] <= 3'b101;
      // memory_array[22009] <= 3'b000;
      // memory_array[22010] <= 3'b000;
      // memory_array[22011] <= 3'b000;
      // memory_array[22012] <= 3'b000;
      // memory_array[22013] <= 3'b000;
      // memory_array[22014] <= 3'b000;
      // memory_array[22015] <= 3'b000;
      // memory_array[22016] <= 3'b000;
      // memory_array[22017] <= 3'b000;
      // memory_array[22018] <= 3'b000;
      // memory_array[22019] <= 3'b000;
      // memory_array[22020] <= 3'b000;
      // memory_array[22021] <= 3'b000;
      // memory_array[22022] <= 3'b000;
      // memory_array[22023] <= 3'b000;
      // memory_array[22024] <= 3'b111;
      // memory_array[22025] <= 3'b111;
      // memory_array[22026] <= 3'b111;
      // memory_array[22027] <= 3'b000;
      // memory_array[22028] <= 3'b000;
      // memory_array[22029] <= 3'b000;
      // memory_array[22030] <= 3'b000;
      // memory_array[22031] <= 3'b000;
      // memory_array[22032] <= 3'b000;
      // memory_array[22033] <= 3'b000;
      // memory_array[22034] <= 3'b000;
      // memory_array[22035] <= 3'b000;
      // memory_array[22036] <= 3'b000;
      // memory_array[22037] <= 3'b111;
      // memory_array[22038] <= 3'b111;
      // memory_array[22039] <= 3'b111;
      // memory_array[22040] <= 3'b111;
      // memory_array[22041] <= 3'b000;
      // memory_array[22042] <= 3'b000;
      // memory_array[22043] <= 3'b111;
      // memory_array[22044] <= 3'b111;
      // memory_array[22045] <= 3'b111;
      // memory_array[22046] <= 3'b111;
      // memory_array[22047] <= 3'b000;
      // memory_array[22048] <= 3'b111;
      // memory_array[22049] <= 3'b101;
      // memory_array[22050] <= 3'b000;
      // memory_array[22051] <= 3'b111;
      // memory_array[22052] <= 3'b111;
      // memory_array[22053] <= 3'b111;
      // memory_array[22054] <= 3'b111;
      // memory_array[22055] <= 3'b000;
      // memory_array[22056] <= 3'b000;
      // memory_array[22057] <= 3'b111;
      // memory_array[22058] <= 3'b111;
      // memory_array[22059] <= 3'b111;
      // memory_array[22060] <= 3'b111;
      // memory_array[22061] <= 3'b000;
      // memory_array[22062] <= 3'b000;
      // memory_array[22063] <= 3'b000;
      // memory_array[22064] <= 3'b000;
      // memory_array[22065] <= 3'b000;
      // memory_array[22066] <= 3'b000;
      // memory_array[22067] <= 3'b111;
      // memory_array[22068] <= 3'b111;
      // memory_array[22069] <= 3'b111;
      // memory_array[22070] <= 3'b111;
      // memory_array[22071] <= 3'b111;
      // memory_array[22072] <= 3'b000;
      // memory_array[22073] <= 3'b000;
      // memory_array[22074] <= 3'b101;
      // memory_array[22075] <= 3'b000;
      // memory_array[22076] <= 3'b000;
      // memory_array[22077] <= 3'b000;
      // memory_array[22078] <= 3'b101;
      // memory_array[22079] <= 3'b101;
      // memory_array[22080] <= 3'b000;
      // memory_array[22081] <= 3'b101;
      // memory_array[22082] <= 3'b000;
      // memory_array[22083] <= 3'b000;
      // memory_array[22084] <= 3'b101;
      // memory_array[22085] <= 3'b000;
      // memory_array[22086] <= 3'b000;
      // memory_array[22087] <= 3'b000;
      // memory_array[22088] <= 3'b000;
      // memory_array[22089] <= 3'b000;
      // memory_array[22090] <= 3'b000;
      // memory_array[22091] <= 3'b111;
      // memory_array[22092] <= 3'b111;
      // memory_array[22093] <= 3'b111;
      // memory_array[22094] <= 3'b111;
      // memory_array[22095] <= 3'b111;
      // memory_array[22096] <= 3'b111;
      // memory_array[22097] <= 3'b111;
      // memory_array[22098] <= 3'b111;
      // memory_array[22099] <= 3'b000;
      // memory_array[22100] <= 3'b000;
      // memory_array[22101] <= 3'b000;
      // memory_array[22102] <= 3'b000;
      // memory_array[22103] <= 3'b000;
      // memory_array[22104] <= 3'b000;
      // memory_array[22105] <= 3'b000;
      // memory_array[22106] <= 3'b000;
      // memory_array[22107] <= 3'b111;
      // memory_array[22108] <= 3'b000;
      // memory_array[22109] <= 3'b000;
      // memory_array[22110] <= 3'b000;
      // memory_array[22111] <= 3'b000;
      // memory_array[22112] <= 3'b000;
      // memory_array[22113] <= 3'b101;
      // memory_array[22114] <= 3'b101;
      // memory_array[22115] <= 3'b000;
      // memory_array[22116] <= 3'b000;
      // memory_array[22117] <= 3'b000;
      // memory_array[22118] <= 3'b000;
      // memory_array[22119] <= 3'b000;
      // memory_array[22120] <= 3'b000;
      // memory_array[22121] <= 3'b000;
      // memory_array[22122] <= 3'b000;
      // memory_array[22123] <= 3'b101;
      // memory_array[22124] <= 3'b000;
      // memory_array[22125] <= 3'b000;
      // memory_array[22126] <= 3'b000;
      // memory_array[22127] <= 3'b000;
      // memory_array[22128] <= 3'b101;
      // memory_array[22129] <= 3'b101;
      // memory_array[22130] <= 3'b000;
      // memory_array[22131] <= 3'b000;
      // memory_array[22132] <= 3'b000;
      // memory_array[22133] <= 3'b000;
      // memory_array[22134] <= 3'b111;
      // memory_array[22135] <= 3'b111;
      // memory_array[22136] <= 3'b111;
      // memory_array[22137] <= 3'b111;
      // memory_array[22138] <= 3'b111;
      // memory_array[22139] <= 3'b000;
      // memory_array[22140] <= 3'b000;
      // memory_array[22141] <= 3'b000;
      // memory_array[22142] <= 3'b111;
      // memory_array[22143] <= 3'b111;
      // memory_array[22144] <= 3'b111;
      // memory_array[22145] <= 3'b111;
      // memory_array[22146] <= 3'b111;
      // memory_array[22147] <= 3'b000;
      // memory_array[22148] <= 3'b111;
      // memory_array[22149] <= 3'b111;
      // memory_array[22150] <= 3'b111;
      // memory_array[22151] <= 3'b111;
      // memory_array[22152] <= 3'b111;
      // memory_array[22153] <= 3'b111;
      // memory_array[22154] <= 3'b111;
      // memory_array[22155] <= 3'b101;
      // memory_array[22156] <= 3'b111;
      // memory_array[22157] <= 3'b111;
      // memory_array[22158] <= 3'b111;
      // memory_array[22159] <= 3'b111;
      // memory_array[22160] <= 3'b000;
      // memory_array[22161] <= 3'b000;
      // memory_array[22162] <= 3'b111;
      // memory_array[22163] <= 3'b111;
      // memory_array[22164] <= 3'b111;
      // memory_array[22165] <= 3'b111;
      // memory_array[22166] <= 3'b111;
      // memory_array[22167] <= 3'b111;
      // memory_array[22168] <= 3'b111;
      // memory_array[22169] <= 3'b111;
      // memory_array[22170] <= 3'b111;
      // memory_array[22171] <= 3'b000;
      // memory_array[22172] <= 3'b000;
      // memory_array[22173] <= 3'b000;
      // memory_array[22174] <= 3'b000;
      // memory_array[22175] <= 3'b111;
      // memory_array[22176] <= 3'b111;
      // memory_array[22177] <= 3'b111;
      // memory_array[22178] <= 3'b111;
      // memory_array[22179] <= 3'b000;
      // memory_array[22180] <= 3'b000;
      // memory_array[22181] <= 3'b000;
      // memory_array[22182] <= 3'b000;
      // memory_array[22183] <= 3'b000;
      // memory_array[22184] <= 3'b000;
      // memory_array[22185] <= 3'b000;
      // memory_array[22186] <= 3'b000;
      // memory_array[22187] <= 3'b000;
      // memory_array[22188] <= 3'b000;
      // memory_array[22189] <= 3'b000;
      // memory_array[22190] <= 3'b000;
      // memory_array[22191] <= 3'b101;
      // memory_array[22192] <= 3'b101;
      // memory_array[22193] <= 3'b110;
      // memory_array[22194] <= 3'b110;
      // memory_array[22195] <= 3'b000;
      // memory_array[22196] <= 3'b000;
      // memory_array[22197] <= 3'b000;
      // memory_array[22198] <= 3'b110;
      // memory_array[22199] <= 3'b101;
      // memory_array[22200] <= 3'b101;
      // memory_array[22201] <= 3'b101;
      // memory_array[22202] <= 3'b101;
      // memory_array[22203] <= 3'b111;
      // memory_array[22204] <= 3'b111;
      // memory_array[22205] <= 3'b101;
      // memory_array[22206] <= 3'b101;
      // memory_array[22207] <= 3'b101;
      // memory_array[22208] <= 3'b101;
      // memory_array[22209] <= 3'b000;
      // memory_array[22210] <= 3'b000;
      // memory_array[22211] <= 3'b110;
      // memory_array[22212] <= 3'b111;
      // memory_array[22213] <= 3'b110;
      // memory_array[22214] <= 3'b110;
      // memory_array[22215] <= 3'b110;
      // memory_array[22216] <= 3'b110;
      // memory_array[22217] <= 3'b111;
      // memory_array[22218] <= 3'b110;
      // memory_array[22219] <= 3'b110;
      // memory_array[22220] <= 3'b111;
      // memory_array[22221] <= 3'b000;
      // memory_array[22222] <= 3'b110;
      // memory_array[22223] <= 3'b000;
      // memory_array[22224] <= 3'b111;
      // memory_array[22225] <= 3'b111;
      // memory_array[22226] <= 3'b111;
      // memory_array[22227] <= 3'b000;
      // memory_array[22228] <= 3'b110;
      // memory_array[22229] <= 3'b110;
      // memory_array[22230] <= 3'b111;
      // memory_array[22231] <= 3'b111;
      // memory_array[22232] <= 3'b000;
      // memory_array[22233] <= 3'b110;
      // memory_array[22234] <= 3'b110;
      // memory_array[22235] <= 3'b110;
      // memory_array[22236] <= 3'b110;
      // memory_array[22237] <= 3'b111;
      // memory_array[22238] <= 3'b111;
      // memory_array[22239] <= 3'b111;
      // memory_array[22240] <= 3'b111;
      // memory_array[22241] <= 3'b000;
      // memory_array[22242] <= 3'b000;
      // memory_array[22243] <= 3'b000;
      // memory_array[22244] <= 3'b111;
      // memory_array[22245] <= 3'b111;
      // memory_array[22246] <= 3'b111;
      // memory_array[22247] <= 3'b111;
      // memory_array[22248] <= 3'b000;
      // memory_array[22249] <= 3'b101;
      // memory_array[22250] <= 3'b000;
      // memory_array[22251] <= 3'b111;
      // memory_array[22252] <= 3'b111;
      // memory_array[22253] <= 3'b111;
      // memory_array[22254] <= 3'b111;
      // memory_array[22255] <= 3'b000;
      // memory_array[22256] <= 3'b000;
      // memory_array[22257] <= 3'b111;
      // memory_array[22258] <= 3'b111;
      // memory_array[22259] <= 3'b111;
      // memory_array[22260] <= 3'b111;
      // memory_array[22261] <= 3'b111;
      // memory_array[22262] <= 3'b111;
      // memory_array[22263] <= 3'b000;
      // memory_array[22264] <= 3'b000;
      // memory_array[22265] <= 3'b000;
      // memory_array[22266] <= 3'b000;
      // memory_array[22267] <= 3'b000;
      // memory_array[22268] <= 3'b000;
      // memory_array[22269] <= 3'b000;
      // memory_array[22270] <= 3'b000;
      // memory_array[22271] <= 3'b000;
      // memory_array[22272] <= 3'b000;
      // memory_array[22273] <= 3'b101;
      // memory_array[22274] <= 3'b101;
      // memory_array[22275] <= 3'b000;
      // memory_array[22276] <= 3'b101;
      // memory_array[22277] <= 3'b101;
      // memory_array[22278] <= 3'b101;
      // memory_array[22279] <= 3'b101;
      // memory_array[22280] <= 3'b000;
      // memory_array[22281] <= 3'b000;
      // memory_array[22282] <= 3'b000;
      // memory_array[22283] <= 3'b101;
      // memory_array[22284] <= 3'b101;
      // memory_array[22285] <= 3'b000;
      // memory_array[22286] <= 3'b000;
      // memory_array[22287] <= 3'b000;
      // memory_array[22288] <= 3'b000;
      // memory_array[22289] <= 3'b101;
      // memory_array[22290] <= 3'b000;
      // memory_array[22291] <= 3'b000;
      // memory_array[22292] <= 3'b000;
      // memory_array[22293] <= 3'b000;
      // memory_array[22294] <= 3'b000;
      // memory_array[22295] <= 3'b000;
      // memory_array[22296] <= 3'b000;
      // memory_array[22297] <= 3'b000;
      // memory_array[22298] <= 3'b000;
      // memory_array[22299] <= 3'b101;
      // memory_array[22300] <= 3'b000;
      // memory_array[22301] <= 3'b101;
      // memory_array[22302] <= 3'b000;
      // memory_array[22303] <= 3'b101;
      // memory_array[22304] <= 3'b000;
      // memory_array[22305] <= 3'b000;
      // memory_array[22306] <= 3'b000;
      // memory_array[22307] <= 3'b000;
      // memory_array[22308] <= 3'b000;
      // memory_array[22309] <= 3'b101;
      // memory_array[22310] <= 3'b000;
      // memory_array[22311] <= 3'b000;
      // memory_array[22312] <= 3'b101;
      // memory_array[22313] <= 3'b000;
      // memory_array[22314] <= 3'b101;
      // memory_array[22315] <= 3'b000;
      // memory_array[22316] <= 3'b101;
      // memory_array[22317] <= 3'b000;
      // memory_array[22318] <= 3'b000;
      // memory_array[22319] <= 3'b000;
      // memory_array[22320] <= 3'b000;
      // memory_array[22321] <= 3'b000;
      // memory_array[22322] <= 3'b000;
      // memory_array[22323] <= 3'b101;
      // memory_array[22324] <= 3'b101;
      // memory_array[22325] <= 3'b000;
      // memory_array[22326] <= 3'b000;
      // memory_array[22327] <= 3'b000;
      // memory_array[22328] <= 3'b101;
      // memory_array[22329] <= 3'b110;
      // memory_array[22330] <= 3'b000;
      // memory_array[22331] <= 3'b000;
      // memory_array[22332] <= 3'b000;
      // memory_array[22333] <= 3'b000;
      // memory_array[22334] <= 3'b000;
      // memory_array[22335] <= 3'b111;
      // memory_array[22336] <= 3'b111;
      // memory_array[22337] <= 3'b111;
      // memory_array[22338] <= 3'b111;
      // memory_array[22339] <= 3'b000;
      // memory_array[22340] <= 3'b000;
      // memory_array[22341] <= 3'b000;
      // memory_array[22342] <= 3'b111;
      // memory_array[22343] <= 3'b111;
      // memory_array[22344] <= 3'b111;
      // memory_array[22345] <= 3'b111;
      // memory_array[22346] <= 3'b111;
      // memory_array[22347] <= 3'b000;
      // memory_array[22348] <= 3'b111;
      // memory_array[22349] <= 3'b111;
      // memory_array[22350] <= 3'b111;
      // memory_array[22351] <= 3'b111;
      // memory_array[22352] <= 3'b111;
      // memory_array[22353] <= 3'b111;
      // memory_array[22354] <= 3'b000;
      // memory_array[22355] <= 3'b000;
      // memory_array[22356] <= 3'b111;
      // memory_array[22357] <= 3'b111;
      // memory_array[22358] <= 3'b111;
      // memory_array[22359] <= 3'b000;
      // memory_array[22360] <= 3'b000;
      // memory_array[22361] <= 3'b000;
      // memory_array[22362] <= 3'b111;
      // memory_array[22363] <= 3'b111;
      // memory_array[22364] <= 3'b111;
      // memory_array[22365] <= 3'b111;
      // memory_array[22366] <= 3'b111;
      // memory_array[22367] <= 3'b111;
      // memory_array[22368] <= 3'b111;
      // memory_array[22369] <= 3'b111;
      // memory_array[22370] <= 3'b111;
      // memory_array[22371] <= 3'b110;
      // memory_array[22372] <= 3'b000;
      // memory_array[22373] <= 3'b110;
      // memory_array[22374] <= 3'b000;
      // memory_array[22375] <= 3'b111;
      // memory_array[22376] <= 3'b111;
      // memory_array[22377] <= 3'b111;
      // memory_array[22378] <= 3'b111;
      // memory_array[22379] <= 3'b110;
      // memory_array[22380] <= 3'b110;
      // memory_array[22381] <= 3'b110;
      // memory_array[22382] <= 3'b110;
      // memory_array[22383] <= 3'b110;
      // memory_array[22384] <= 3'b110;
      // memory_array[22385] <= 3'b111;
      // memory_array[22386] <= 3'b111;
      // memory_array[22387] <= 3'b111;
      // memory_array[22388] <= 3'b110;
      // memory_array[22389] <= 3'b000;
      // memory_array[22390] <= 3'b000;
      // memory_array[22391] <= 3'b101;
      // memory_array[22392] <= 3'b101;
      // memory_array[22393] <= 3'b101;
      // memory_array[22394] <= 3'b101;
      // memory_array[22395] <= 3'b111;
      // memory_array[22396] <= 3'b111;
      // memory_array[22397] <= 3'b101;
      // memory_array[22398] <= 3'b101;
      // memory_array[22399] <= 3'b101;
      // memory_array[22400] <= 3'b101;
      // memory_array[22401] <= 3'b101;
      // memory_array[22402] <= 3'b101;
      // memory_array[22403] <= 3'b101;
      // memory_array[22404] <= 3'b101;
      // memory_array[22405] <= 3'b101;
      // memory_array[22406] <= 3'b101;
      // memory_array[22407] <= 3'b101;
      // memory_array[22408] <= 3'b101;
      // memory_array[22409] <= 3'b000;
      // memory_array[22410] <= 3'b000;
      // memory_array[22411] <= 3'b110;
      // memory_array[22412] <= 3'b111;
      // memory_array[22413] <= 3'b110;
      // memory_array[22414] <= 3'b110;
      // memory_array[22415] <= 3'b110;
      // memory_array[22416] <= 3'b110;
      // memory_array[22417] <= 3'b111;
      // memory_array[22418] <= 3'b110;
      // memory_array[22419] <= 3'b110;
      // memory_array[22420] <= 3'b111;
      // memory_array[22421] <= 3'b000;
      // memory_array[22422] <= 3'b110;
      // memory_array[22423] <= 3'b000;
      // memory_array[22424] <= 3'b111;
      // memory_array[22425] <= 3'b111;
      // memory_array[22426] <= 3'b111;
      // memory_array[22427] <= 3'b000;
      // memory_array[22428] <= 3'b110;
      // memory_array[22429] <= 3'b110;
      // memory_array[22430] <= 3'b111;
      // memory_array[22431] <= 3'b111;
      // memory_array[22432] <= 3'b000;
      // memory_array[22433] <= 3'b110;
      // memory_array[22434] <= 3'b110;
      // memory_array[22435] <= 3'b110;
      // memory_array[22436] <= 3'b110;
      // memory_array[22437] <= 3'b111;
      // memory_array[22438] <= 3'b111;
      // memory_array[22439] <= 3'b111;
      // memory_array[22440] <= 3'b111;
      // memory_array[22441] <= 3'b000;
      // memory_array[22442] <= 3'b000;
      // memory_array[22443] <= 3'b110;
      // memory_array[22444] <= 3'b111;
      // memory_array[22445] <= 3'b111;
      // memory_array[22446] <= 3'b111;
      // memory_array[22447] <= 3'b111;
      // memory_array[22448] <= 3'b111;
      // memory_array[22449] <= 3'b000;
      // memory_array[22450] <= 3'b000;
      // memory_array[22451] <= 3'b111;
      // memory_array[22452] <= 3'b111;
      // memory_array[22453] <= 3'b111;
      // memory_array[22454] <= 3'b111;
      // memory_array[22455] <= 3'b111;
      // memory_array[22456] <= 3'b111;
      // memory_array[22457] <= 3'b111;
      // memory_array[22458] <= 3'b111;
      // memory_array[22459] <= 3'b000;
      // memory_array[22460] <= 3'b000;
      // memory_array[22461] <= 3'b000;
      // memory_array[22462] <= 3'b000;
      // memory_array[22463] <= 3'b000;
      // memory_array[22464] <= 3'b000;
      // memory_array[22465] <= 3'b000;
      // memory_array[22466] <= 3'b000;
      // memory_array[22467] <= 3'b000;
      // memory_array[22468] <= 3'b101;
      // memory_array[22469] <= 3'b000;
      // memory_array[22470] <= 3'b000;
      // memory_array[22471] <= 3'b000;
      // memory_array[22472] <= 3'b000;
      // memory_array[22473] <= 3'b101;
      // memory_array[22474] <= 3'b101;
      // memory_array[22475] <= 3'b000;
      // memory_array[22476] <= 3'b000;
      // memory_array[22477] <= 3'b000;
      // memory_array[22478] <= 3'b101;
      // memory_array[22479] <= 3'b101;
      // memory_array[22480] <= 3'b000;
      // memory_array[22481] <= 3'b000;
      // memory_array[22482] <= 3'b000;
      // memory_array[22483] <= 3'b000;
      // memory_array[22484] <= 3'b000;
      // memory_array[22485] <= 3'b000;
      // memory_array[22486] <= 3'b000;
      // memory_array[22487] <= 3'b000;
      // memory_array[22488] <= 3'b101;
      // memory_array[22489] <= 3'b101;
      // memory_array[22490] <= 3'b000;
      // memory_array[22491] <= 3'b000;
      // memory_array[22492] <= 3'b000;
      // memory_array[22493] <= 3'b101;
      // memory_array[22494] <= 3'b101;
      // memory_array[22495] <= 3'b000;
      // memory_array[22496] <= 3'b000;
      // memory_array[22497] <= 3'b000;
      // memory_array[22498] <= 3'b110;
      // memory_array[22499] <= 3'b000;
      // memory_array[22500] <= 3'b000;
      // memory_array[22501] <= 3'b000;
      // memory_array[22502] <= 3'b000;
      // memory_array[22503] <= 3'b000;
      // memory_array[22504] <= 3'b101;
      // memory_array[22505] <= 3'b000;
      // memory_array[22506] <= 3'b101;
      // memory_array[22507] <= 3'b101;
      // memory_array[22508] <= 3'b000;
      // memory_array[22509] <= 3'b101;
      // memory_array[22510] <= 3'b101;
      // memory_array[22511] <= 3'b000;
      // memory_array[22512] <= 3'b000;
      // memory_array[22513] <= 3'b000;
      // memory_array[22514] <= 3'b000;
      // memory_array[22515] <= 3'b000;
      // memory_array[22516] <= 3'b000;
      // memory_array[22517] <= 3'b000;
      // memory_array[22518] <= 3'b000;
      // memory_array[22519] <= 3'b000;
      // memory_array[22520] <= 3'b000;
      // memory_array[22521] <= 3'b000;
      // memory_array[22522] <= 3'b000;
      // memory_array[22523] <= 3'b101;
      // memory_array[22524] <= 3'b101;
      // memory_array[22525] <= 3'b000;
      // memory_array[22526] <= 3'b000;
      // memory_array[22527] <= 3'b000;
      // memory_array[22528] <= 3'b101;
      // memory_array[22529] <= 3'b101;
      // memory_array[22530] <= 3'b000;
      // memory_array[22531] <= 3'b000;
      // memory_array[22532] <= 3'b000;
      // memory_array[22533] <= 3'b000;
      // memory_array[22534] <= 3'b000;
      // memory_array[22535] <= 3'b000;
      // memory_array[22536] <= 3'b000;
      // memory_array[22537] <= 3'b000;
      // memory_array[22538] <= 3'b101;
      // memory_array[22539] <= 3'b000;
      // memory_array[22540] <= 3'b000;
      // memory_array[22541] <= 3'b000;
      // memory_array[22542] <= 3'b111;
      // memory_array[22543] <= 3'b111;
      // memory_array[22544] <= 3'b111;
      // memory_array[22545] <= 3'b111;
      // memory_array[22546] <= 3'b111;
      // memory_array[22547] <= 3'b111;
      // memory_array[22548] <= 3'b000;
      // memory_array[22549] <= 3'b111;
      // memory_array[22550] <= 3'b111;
      // memory_array[22551] <= 3'b111;
      // memory_array[22552] <= 3'b111;
      // memory_array[22553] <= 3'b111;
      // memory_array[22554] <= 3'b111;
      // memory_array[22555] <= 3'b111;
      // memory_array[22556] <= 3'b111;
      // memory_array[22557] <= 3'b111;
      // memory_array[22558] <= 3'b000;
      // memory_array[22559] <= 3'b110;
      // memory_array[22560] <= 3'b000;
      // memory_array[22561] <= 3'b000;
      // memory_array[22562] <= 3'b111;
      // memory_array[22563] <= 3'b111;
      // memory_array[22564] <= 3'b111;
      // memory_array[22565] <= 3'b111;
      // memory_array[22566] <= 3'b111;
      // memory_array[22567] <= 3'b111;
      // memory_array[22568] <= 3'b111;
      // memory_array[22569] <= 3'b111;
      // memory_array[22570] <= 3'b111;
      // memory_array[22571] <= 3'b000;
      // memory_array[22572] <= 3'b000;
      // memory_array[22573] <= 3'b110;
      // memory_array[22574] <= 3'b000;
      // memory_array[22575] <= 3'b111;
      // memory_array[22576] <= 3'b111;
      // memory_array[22577] <= 3'b111;
      // memory_array[22578] <= 3'b111;
      // memory_array[22579] <= 3'b110;
      // memory_array[22580] <= 3'b110;
      // memory_array[22581] <= 3'b110;
      // memory_array[22582] <= 3'b110;
      // memory_array[22583] <= 3'b110;
      // memory_array[22584] <= 3'b110;
      // memory_array[22585] <= 3'b111;
      // memory_array[22586] <= 3'b111;
      // memory_array[22587] <= 3'b111;
      // memory_array[22588] <= 3'b110;
      // memory_array[22589] <= 3'b000;
      // memory_array[22590] <= 3'b000;
      // memory_array[22591] <= 3'b101;
      // memory_array[22592] <= 3'b111;
      // memory_array[22593] <= 3'b101;
      // memory_array[22594] <= 3'b101;
      // memory_array[22595] <= 3'b101;
      // memory_array[22596] <= 3'b101;
      // memory_array[22597] <= 3'b101;
      // memory_array[22598] <= 3'b101;
      // memory_array[22599] <= 3'b101;
      // memory_array[22600] <= 3'b101;
      // memory_array[22601] <= 3'b101;
      // memory_array[22602] <= 3'b101;
      // memory_array[22603] <= 3'b101;
      // memory_array[22604] <= 3'b101;
      // memory_array[22605] <= 3'b101;
      // memory_array[22606] <= 3'b101;
      // memory_array[22607] <= 3'b101;
      // memory_array[22608] <= 3'b101;
      // memory_array[22609] <= 3'b000;
      // memory_array[22610] <= 3'b000;
      // memory_array[22611] <= 3'b110;
      // memory_array[22612] <= 3'b110;
      // memory_array[22613] <= 3'b111;
      // memory_array[22614] <= 3'b111;
      // memory_array[22615] <= 3'b110;
      // memory_array[22616] <= 3'b110;
      // memory_array[22617] <= 3'b110;
      // memory_array[22618] <= 3'b111;
      // memory_array[22619] <= 3'b111;
      // memory_array[22620] <= 3'b110;
      // memory_array[22621] <= 3'b000;
      // memory_array[22622] <= 3'b110;
      // memory_array[22623] <= 3'b000;
      // memory_array[22624] <= 3'b111;
      // memory_array[22625] <= 3'b111;
      // memory_array[22626] <= 3'b111;
      // memory_array[22627] <= 3'b000;
      // memory_array[22628] <= 3'b111;
      // memory_array[22629] <= 3'b111;
      // memory_array[22630] <= 3'b110;
      // memory_array[22631] <= 3'b110;
      // memory_array[22632] <= 3'b000;
      // memory_array[22633] <= 3'b111;
      // memory_array[22634] <= 3'b110;
      // memory_array[22635] <= 3'b110;
      // memory_array[22636] <= 3'b110;
      // memory_array[22637] <= 3'b111;
      // memory_array[22638] <= 3'b111;
      // memory_array[22639] <= 3'b111;
      // memory_array[22640] <= 3'b111;
      // memory_array[22641] <= 3'b000;
      // memory_array[22642] <= 3'b110;
      // memory_array[22643] <= 3'b000;
      // memory_array[22644] <= 3'b000;
      // memory_array[22645] <= 3'b111;
      // memory_array[22646] <= 3'b111;
      // memory_array[22647] <= 3'b111;
      // memory_array[22648] <= 3'b111;
      // memory_array[22649] <= 3'b111;
      // memory_array[22650] <= 3'b111;
      // memory_array[22651] <= 3'b111;
      // memory_array[22652] <= 3'b111;
      // memory_array[22653] <= 3'b111;
      // memory_array[22654] <= 3'b111;
      // memory_array[22655] <= 3'b111;
      // memory_array[22656] <= 3'b000;
      // memory_array[22657] <= 3'b000;
      // memory_array[22658] <= 3'b000;
      // memory_array[22659] <= 3'b000;
      // memory_array[22660] <= 3'b000;
      // memory_array[22661] <= 3'b000;
      // memory_array[22662] <= 3'b000;
      // memory_array[22663] <= 3'b000;
      // memory_array[22664] <= 3'b000;
      // memory_array[22665] <= 3'b000;
      // memory_array[22666] <= 3'b000;
      // memory_array[22667] <= 3'b000;
      // memory_array[22668] <= 3'b000;
      // memory_array[22669] <= 3'b000;
      // memory_array[22670] <= 3'b101;
      // memory_array[22671] <= 3'b101;
      // memory_array[22672] <= 3'b101;
      // memory_array[22673] <= 3'b000;
      // memory_array[22674] <= 3'b000;
      // memory_array[22675] <= 3'b101;
      // memory_array[22676] <= 3'b101;
      // memory_array[22677] <= 3'b101;
      // memory_array[22678] <= 3'b000;
      // memory_array[22679] <= 3'b000;
      // memory_array[22680] <= 3'b000;
      // memory_array[22681] <= 3'b000;
      // memory_array[22682] <= 3'b000;
      // memory_array[22683] <= 3'b000;
      // memory_array[22684] <= 3'b000;
      // memory_array[22685] <= 3'b000;
      // memory_array[22686] <= 3'b000;
      // memory_array[22687] <= 3'b000;
      // memory_array[22688] <= 3'b000;
      // memory_array[22689] <= 3'b000;
      // memory_array[22690] <= 3'b101;
      // memory_array[22691] <= 3'b101;
      // memory_array[22692] <= 3'b101;
      // memory_array[22693] <= 3'b000;
      // memory_array[22694] <= 3'b000;
      // memory_array[22695] <= 3'b101;
      // memory_array[22696] <= 3'b000;
      // memory_array[22697] <= 3'b110;
      // memory_array[22698] <= 3'b000;
      // memory_array[22699] <= 3'b000;
      // memory_array[22700] <= 3'b000;
      // memory_array[22701] <= 3'b000;
      // memory_array[22702] <= 3'b000;
      // memory_array[22703] <= 3'b000;
      // memory_array[22704] <= 3'b101;
      // memory_array[22705] <= 3'b101;
      // memory_array[22706] <= 3'b000;
      // memory_array[22707] <= 3'b000;
      // memory_array[22708] <= 3'b000;
      // memory_array[22709] <= 3'b101;
      // memory_array[22710] <= 3'b101;
      // memory_array[22711] <= 3'b101;
      // memory_array[22712] <= 3'b101;
      // memory_array[22713] <= 3'b101;
      // memory_array[22714] <= 3'b101;
      // memory_array[22715] <= 3'b000;
      // memory_array[22716] <= 3'b000;
      // memory_array[22717] <= 3'b000;
      // memory_array[22718] <= 3'b101;
      // memory_array[22719] <= 3'b000;
      // memory_array[22720] <= 3'b000;
      // memory_array[22721] <= 3'b101;
      // memory_array[22722] <= 3'b101;
      // memory_array[22723] <= 3'b000;
      // memory_array[22724] <= 3'b000;
      // memory_array[22725] <= 3'b101;
      // memory_array[22726] <= 3'b101;
      // memory_array[22727] <= 3'b000;
      // memory_array[22728] <= 3'b000;
      // memory_array[22729] <= 3'b000;
      // memory_array[22730] <= 3'b000;
      // memory_array[22731] <= 3'b000;
      // memory_array[22732] <= 3'b000;
      // memory_array[22733] <= 3'b000;
      // memory_array[22734] <= 3'b000;
      // memory_array[22735] <= 3'b000;
      // memory_array[22736] <= 3'b000;
      // memory_array[22737] <= 3'b101;
      // memory_array[22738] <= 3'b000;
      // memory_array[22739] <= 3'b000;
      // memory_array[22740] <= 3'b101;
      // memory_array[22741] <= 3'b000;
      // memory_array[22742] <= 3'b000;
      // memory_array[22743] <= 3'b000;
      // memory_array[22744] <= 3'b111;
      // memory_array[22745] <= 3'b111;
      // memory_array[22746] <= 3'b111;
      // memory_array[22747] <= 3'b111;
      // memory_array[22748] <= 3'b111;
      // memory_array[22749] <= 3'b111;
      // memory_array[22750] <= 3'b111;
      // memory_array[22751] <= 3'b111;
      // memory_array[22752] <= 3'b111;
      // memory_array[22753] <= 3'b111;
      // memory_array[22754] <= 3'b111;
      // memory_array[22755] <= 3'b111;
      // memory_array[22756] <= 3'b000;
      // memory_array[22757] <= 3'b000;
      // memory_array[22758] <= 3'b000;
      // memory_array[22759] <= 3'b000;
      // memory_array[22760] <= 3'b110;
      // memory_array[22761] <= 3'b000;
      // memory_array[22762] <= 3'b111;
      // memory_array[22763] <= 3'b111;
      // memory_array[22764] <= 3'b111;
      // memory_array[22765] <= 3'b111;
      // memory_array[22766] <= 3'b000;
      // memory_array[22767] <= 3'b111;
      // memory_array[22768] <= 3'b111;
      // memory_array[22769] <= 3'b111;
      // memory_array[22770] <= 3'b111;
      // memory_array[22771] <= 3'b000;
      // memory_array[22772] <= 3'b000;
      // memory_array[22773] <= 3'b110;
      // memory_array[22774] <= 3'b000;
      // memory_array[22775] <= 3'b111;
      // memory_array[22776] <= 3'b111;
      // memory_array[22777] <= 3'b111;
      // memory_array[22778] <= 3'b111;
      // memory_array[22779] <= 3'b110;
      // memory_array[22780] <= 3'b110;
      // memory_array[22781] <= 3'b110;
      // memory_array[22782] <= 3'b110;
      // memory_array[22783] <= 3'b000;
      // memory_array[22784] <= 3'b110;
      // memory_array[22785] <= 3'b110;
      // memory_array[22786] <= 3'b110;
      // memory_array[22787] <= 3'b110;
      // memory_array[22788] <= 3'b110;
      // memory_array[22789] <= 3'b000;
      // memory_array[22790] <= 3'b000;
      // memory_array[22791] <= 3'b101;
      // memory_array[22792] <= 3'b101;
      // memory_array[22793] <= 3'b101;
      // memory_array[22794] <= 3'b101;
      // memory_array[22795] <= 3'b101;
      // memory_array[22796] <= 3'b101;
      // memory_array[22797] <= 3'b101;
      // memory_array[22798] <= 3'b101;
      // memory_array[22799] <= 3'b101;
      // memory_array[22800] <= 3'b101;
      // memory_array[22801] <= 3'b101;
      // memory_array[22802] <= 3'b101;
      // memory_array[22803] <= 3'b111;
      // memory_array[22804] <= 3'b111;
      // memory_array[22805] <= 3'b101;
      // memory_array[22806] <= 3'b101;
      // memory_array[22807] <= 3'b101;
      // memory_array[22808] <= 3'b101;
      // memory_array[22809] <= 3'b000;
      // memory_array[22810] <= 3'b000;
      // memory_array[22811] <= 3'b110;
      // memory_array[22812] <= 3'b111;
      // memory_array[22813] <= 3'b110;
      // memory_array[22814] <= 3'b110;
      // memory_array[22815] <= 3'b110;
      // memory_array[22816] <= 3'b110;
      // memory_array[22817] <= 3'b111;
      // memory_array[22818] <= 3'b110;
      // memory_array[22819] <= 3'b110;
      // memory_array[22820] <= 3'b111;
      // memory_array[22821] <= 3'b000;
      // memory_array[22822] <= 3'b110;
      // memory_array[22823] <= 3'b000;
      // memory_array[22824] <= 3'b111;
      // memory_array[22825] <= 3'b111;
      // memory_array[22826] <= 3'b111;
      // memory_array[22827] <= 3'b000;
      // memory_array[22828] <= 3'b110;
      // memory_array[22829] <= 3'b110;
      // memory_array[22830] <= 3'b111;
      // memory_array[22831] <= 3'b111;
      // memory_array[22832] <= 3'b000;
      // memory_array[22833] <= 3'b110;
      // memory_array[22834] <= 3'b110;
      // memory_array[22835] <= 3'b110;
      // memory_array[22836] <= 3'b110;
      // memory_array[22837] <= 3'b111;
      // memory_array[22838] <= 3'b111;
      // memory_array[22839] <= 3'b111;
      // memory_array[22840] <= 3'b111;
      // memory_array[22841] <= 3'b000;
      // memory_array[22842] <= 3'b000;
      // memory_array[22843] <= 3'b110;
      // memory_array[22844] <= 3'b000;
      // memory_array[22845] <= 3'b111;
      // memory_array[22846] <= 3'b111;
      // memory_array[22847] <= 3'b111;
      // memory_array[22848] <= 3'b111;
      // memory_array[22849] <= 3'b111;
      // memory_array[22850] <= 3'b111;
      // memory_array[22851] <= 3'b111;
      // memory_array[22852] <= 3'b111;
      // memory_array[22853] <= 3'b111;
      // memory_array[22854] <= 3'b000;
      // memory_array[22855] <= 3'b000;
      // memory_array[22856] <= 3'b000;
      // memory_array[22857] <= 3'b000;
      // memory_array[22858] <= 3'b000;
      // memory_array[22859] <= 3'b000;
      // memory_array[22860] <= 3'b000;
      // memory_array[22861] <= 3'b000;
      // memory_array[22862] <= 3'b000;
      // memory_array[22863] <= 3'b000;
      // memory_array[22864] <= 3'b000;
      // memory_array[22865] <= 3'b000;
      // memory_array[22866] <= 3'b000;
      // memory_array[22867] <= 3'b000;
      // memory_array[22868] <= 3'b101;
      // memory_array[22869] <= 3'b000;
      // memory_array[22870] <= 3'b000;
      // memory_array[22871] <= 3'b000;
      // memory_array[22872] <= 3'b000;
      // memory_array[22873] <= 3'b000;
      // memory_array[22874] <= 3'b000;
      // memory_array[22875] <= 3'b000;
      // memory_array[22876] <= 3'b000;
      // memory_array[22877] <= 3'b000;
      // memory_array[22878] <= 3'b000;
      // memory_array[22879] <= 3'b000;
      // memory_array[22880] <= 3'b000;
      // memory_array[22881] <= 3'b000;
      // memory_array[22882] <= 3'b000;
      // memory_array[22883] <= 3'b000;
      // memory_array[22884] <= 3'b101;
      // memory_array[22885] <= 3'b000;
      // memory_array[22886] <= 3'b000;
      // memory_array[22887] <= 3'b000;
      // memory_array[22888] <= 3'b101;
      // memory_array[22889] <= 3'b101;
      // memory_array[22890] <= 3'b000;
      // memory_array[22891] <= 3'b000;
      // memory_array[22892] <= 3'b000;
      // memory_array[22893] <= 3'b101;
      // memory_array[22894] <= 3'b101;
      // memory_array[22895] <= 3'b000;
      // memory_array[22896] <= 3'b000;
      // memory_array[22897] <= 3'b000;
      // memory_array[22898] <= 3'b000;
      // memory_array[22899] <= 3'b000;
      // memory_array[22900] <= 3'b000;
      // memory_array[22901] <= 3'b000;
      // memory_array[22902] <= 3'b000;
      // memory_array[22903] <= 3'b101;
      // memory_array[22904] <= 3'b000;
      // memory_array[22905] <= 3'b000;
      // memory_array[22906] <= 3'b000;
      // memory_array[22907] <= 3'b000;
      // memory_array[22908] <= 3'b101;
      // memory_array[22909] <= 3'b101;
      // memory_array[22910] <= 3'b101;
      // memory_array[22911] <= 3'b101;
      // memory_array[22912] <= 3'b101;
      // memory_array[22913] <= 3'b101;
      // memory_array[22914] <= 3'b101;
      // memory_array[22915] <= 3'b101;
      // memory_array[22916] <= 3'b101;
      // memory_array[22917] <= 3'b000;
      // memory_array[22918] <= 3'b000;
      // memory_array[22919] <= 3'b000;
      // memory_array[22920] <= 3'b000;
      // memory_array[22921] <= 3'b000;
      // memory_array[22922] <= 3'b000;
      // memory_array[22923] <= 3'b101;
      // memory_array[22924] <= 3'b101;
      // memory_array[22925] <= 3'b000;
      // memory_array[22926] <= 3'b000;
      // memory_array[22927] <= 3'b000;
      // memory_array[22928] <= 3'b101;
      // memory_array[22929] <= 3'b000;
      // memory_array[22930] <= 3'b000;
      // memory_array[22931] <= 3'b000;
      // memory_array[22932] <= 3'b000;
      // memory_array[22933] <= 3'b000;
      // memory_array[22934] <= 3'b000;
      // memory_array[22935] <= 3'b000;
      // memory_array[22936] <= 3'b000;
      // memory_array[22937] <= 3'b000;
      // memory_array[22938] <= 3'b000;
      // memory_array[22939] <= 3'b000;
      // memory_array[22940] <= 3'b000;
      // memory_array[22941] <= 3'b000;
      // memory_array[22942] <= 3'b000;
      // memory_array[22943] <= 3'b000;
      // memory_array[22944] <= 3'b000;
      // memory_array[22945] <= 3'b000;
      // memory_array[22946] <= 3'b000;
      // memory_array[22947] <= 3'b111;
      // memory_array[22948] <= 3'b111;
      // memory_array[22949] <= 3'b111;
      // memory_array[22950] <= 3'b111;
      // memory_array[22951] <= 3'b111;
      // memory_array[22952] <= 3'b111;
      // memory_array[22953] <= 3'b111;
      // memory_array[22954] <= 3'b111;
      // memory_array[22955] <= 3'b000;
      // memory_array[22956] <= 3'b110;
      // memory_array[22957] <= 3'b000;
      // memory_array[22958] <= 3'b110;
      // memory_array[22959] <= 3'b110;
      // memory_array[22960] <= 3'b000;
      // memory_array[22961] <= 3'b000;
      // memory_array[22962] <= 3'b111;
      // memory_array[22963] <= 3'b111;
      // memory_array[22964] <= 3'b111;
      // memory_array[22965] <= 3'b111;
      // memory_array[22966] <= 3'b000;
      // memory_array[22967] <= 3'b111;
      // memory_array[22968] <= 3'b111;
      // memory_array[22969] <= 3'b111;
      // memory_array[22970] <= 3'b111;
      // memory_array[22971] <= 3'b000;
      // memory_array[22972] <= 3'b000;
      // memory_array[22973] <= 3'b110;
      // memory_array[22974] <= 3'b000;
      // memory_array[22975] <= 3'b111;
      // memory_array[22976] <= 3'b111;
      // memory_array[22977] <= 3'b111;
      // memory_array[22978] <= 3'b111;
      // memory_array[22979] <= 3'b110;
      // memory_array[22980] <= 3'b110;
      // memory_array[22981] <= 3'b110;
      // memory_array[22982] <= 3'b110;
      // memory_array[22983] <= 3'b110;
      // memory_array[22984] <= 3'b110;
      // memory_array[22985] <= 3'b111;
      // memory_array[22986] <= 3'b111;
      // memory_array[22987] <= 3'b111;
      // memory_array[22988] <= 3'b110;
      // memory_array[22989] <= 3'b000;
      // memory_array[22990] <= 3'b000;
      // memory_array[22991] <= 3'b101;
      // memory_array[22992] <= 3'b101;
      // memory_array[22993] <= 3'b101;
      // memory_array[22994] <= 3'b101;
      // memory_array[22995] <= 3'b111;
      // memory_array[22996] <= 3'b111;
      // memory_array[22997] <= 3'b101;
      // memory_array[22998] <= 3'b101;
      // memory_array[22999] <= 3'b101;
      // memory_array[23000] <= 3'b101;
      // memory_array[23001] <= 3'b101;
      // memory_array[23002] <= 3'b110;
      // memory_array[23003] <= 3'b101;
      // memory_array[23004] <= 3'b101;
      // memory_array[23005] <= 3'b110;
      // memory_array[23006] <= 3'b101;
      // memory_array[23007] <= 3'b101;
      // memory_array[23008] <= 3'b101;
      // memory_array[23009] <= 3'b000;
      // memory_array[23010] <= 3'b000;
      // memory_array[23011] <= 3'b110;
      // memory_array[23012] <= 3'b110;
      // memory_array[23013] <= 3'b110;
      // memory_array[23014] <= 3'b110;
      // memory_array[23015] <= 3'b110;
      // memory_array[23016] <= 3'b110;
      // memory_array[23017] <= 3'b110;
      // memory_array[23018] <= 3'b110;
      // memory_array[23019] <= 3'b110;
      // memory_array[23020] <= 3'b110;
      // memory_array[23021] <= 3'b000;
      // memory_array[23022] <= 3'b110;
      // memory_array[23023] <= 3'b000;
      // memory_array[23024] <= 3'b111;
      // memory_array[23025] <= 3'b111;
      // memory_array[23026] <= 3'b111;
      // memory_array[23027] <= 3'b000;
      // memory_array[23028] <= 3'b111;
      // memory_array[23029] <= 3'b110;
      // memory_array[23030] <= 3'b110;
      // memory_array[23031] <= 3'b110;
      // memory_array[23032] <= 3'b000;
      // memory_array[23033] <= 3'b110;
      // memory_array[23034] <= 3'b000;
      // memory_array[23035] <= 3'b110;
      // memory_array[23036] <= 3'b110;
      // memory_array[23037] <= 3'b111;
      // memory_array[23038] <= 3'b111;
      // memory_array[23039] <= 3'b111;
      // memory_array[23040] <= 3'b111;
      // memory_array[23041] <= 3'b000;
      // memory_array[23042] <= 3'b110;
      // memory_array[23043] <= 3'b000;
      // memory_array[23044] <= 3'b111;
      // memory_array[23045] <= 3'b000;
      // memory_array[23046] <= 3'b111;
      // memory_array[23047] <= 3'b111;
      // memory_array[23048] <= 3'b111;
      // memory_array[23049] <= 3'b111;
      // memory_array[23050] <= 3'b111;
      // memory_array[23051] <= 3'b000;
      // memory_array[23052] <= 3'b000;
      // memory_array[23053] <= 3'b000;
      // memory_array[23054] <= 3'b000;
      // memory_array[23055] <= 3'b000;
      // memory_array[23056] <= 3'b000;
      // memory_array[23057] <= 3'b000;
      // memory_array[23058] <= 3'b000;
      // memory_array[23059] <= 3'b000;
      // memory_array[23060] <= 3'b000;
      // memory_array[23061] <= 3'b000;
      // memory_array[23062] <= 3'b000;
      // memory_array[23063] <= 3'b000;
      // memory_array[23064] <= 3'b000;
      // memory_array[23065] <= 3'b000;
      // memory_array[23066] <= 3'b101;
      // memory_array[23067] <= 3'b101;
      // memory_array[23068] <= 3'b000;
      // memory_array[23069] <= 3'b000;
      // memory_array[23070] <= 3'b000;
      // memory_array[23071] <= 3'b000;
      // memory_array[23072] <= 3'b000;
      // memory_array[23073] <= 3'b000;
      // memory_array[23074] <= 3'b000;
      // memory_array[23075] <= 3'b000;
      // memory_array[23076] <= 3'b000;
      // memory_array[23077] <= 3'b000;
      // memory_array[23078] <= 3'b000;
      // memory_array[23079] <= 3'b000;
      // memory_array[23080] <= 3'b000;
      // memory_array[23081] <= 3'b000;
      // memory_array[23082] <= 3'b000;
      // memory_array[23083] <= 3'b000;
      // memory_array[23084] <= 3'b000;
      // memory_array[23085] <= 3'b000;
      // memory_array[23086] <= 3'b000;
      // memory_array[23087] <= 3'b000;
      // memory_array[23088] <= 3'b000;
      // memory_array[23089] <= 3'b000;
      // memory_array[23090] <= 3'b101;
      // memory_array[23091] <= 3'b101;
      // memory_array[23092] <= 3'b101;
      // memory_array[23093] <= 3'b000;
      // memory_array[23094] <= 3'b000;
      // memory_array[23095] <= 3'b000;
      // memory_array[23096] <= 3'b110;
      // memory_array[23097] <= 3'b000;
      // memory_array[23098] <= 3'b000;
      // memory_array[23099] <= 3'b000;
      // memory_array[23100] <= 3'b000;
      // memory_array[23101] <= 3'b101;
      // memory_array[23102] <= 3'b000;
      // memory_array[23103] <= 3'b000;
      // memory_array[23104] <= 3'b000;
      // memory_array[23105] <= 3'b000;
      // memory_array[23106] <= 3'b000;
      // memory_array[23107] <= 3'b000;
      // memory_array[23108] <= 3'b000;
      // memory_array[23109] <= 3'b101;
      // memory_array[23110] <= 3'b101;
      // memory_array[23111] <= 3'b101;
      // memory_array[23112] <= 3'b101;
      // memory_array[23113] <= 3'b101;
      // memory_array[23114] <= 3'b101;
      // memory_array[23115] <= 3'b101;
      // memory_array[23116] <= 3'b101;
      // memory_array[23117] <= 3'b101;
      // memory_array[23118] <= 3'b000;
      // memory_array[23119] <= 3'b000;
      // memory_array[23120] <= 3'b000;
      // memory_array[23121] <= 3'b000;
      // memory_array[23122] <= 3'b101;
      // memory_array[23123] <= 3'b000;
      // memory_array[23124] <= 3'b000;
      // memory_array[23125] <= 3'b101;
      // memory_array[23126] <= 3'b101;
      // memory_array[23127] <= 3'b101;
      // memory_array[23128] <= 3'b000;
      // memory_array[23129] <= 3'b000;
      // memory_array[23130] <= 3'b000;
      // memory_array[23131] <= 3'b000;
      // memory_array[23132] <= 3'b000;
      // memory_array[23133] <= 3'b000;
      // memory_array[23134] <= 3'b000;
      // memory_array[23135] <= 3'b000;
      // memory_array[23136] <= 3'b000;
      // memory_array[23137] <= 3'b000;
      // memory_array[23138] <= 3'b000;
      // memory_array[23139] <= 3'b000;
      // memory_array[23140] <= 3'b000;
      // memory_array[23141] <= 3'b000;
      // memory_array[23142] <= 3'b000;
      // memory_array[23143] <= 3'b000;
      // memory_array[23144] <= 3'b000;
      // memory_array[23145] <= 3'b000;
      // memory_array[23146] <= 3'b000;
      // memory_array[23147] <= 3'b000;
      // memory_array[23148] <= 3'b000;
      // memory_array[23149] <= 3'b000;
      // memory_array[23150] <= 3'b111;
      // memory_array[23151] <= 3'b111;
      // memory_array[23152] <= 3'b111;
      // memory_array[23153] <= 3'b111;
      // memory_array[23154] <= 3'b000;
      // memory_array[23155] <= 3'b101;
      // memory_array[23156] <= 3'b110;
      // memory_array[23157] <= 3'b110;
      // memory_array[23158] <= 3'b000;
      // memory_array[23159] <= 3'b000;
      // memory_array[23160] <= 3'b110;
      // memory_array[23161] <= 3'b000;
      // memory_array[23162] <= 3'b111;
      // memory_array[23163] <= 3'b111;
      // memory_array[23164] <= 3'b111;
      // memory_array[23165] <= 3'b111;
      // memory_array[23166] <= 3'b000;
      // memory_array[23167] <= 3'b111;
      // memory_array[23168] <= 3'b111;
      // memory_array[23169] <= 3'b111;
      // memory_array[23170] <= 3'b111;
      // memory_array[23171] <= 3'b111;
      // memory_array[23172] <= 3'b000;
      // memory_array[23173] <= 3'b111;
      // memory_array[23174] <= 3'b000;
      // memory_array[23175] <= 3'b111;
      // memory_array[23176] <= 3'b111;
      // memory_array[23177] <= 3'b111;
      // memory_array[23178] <= 3'b111;
      // memory_array[23179] <= 3'b110;
      // memory_array[23180] <= 3'b110;
      // memory_array[23181] <= 3'b110;
      // memory_array[23182] <= 3'b110;
      // memory_array[23183] <= 3'b000;
      // memory_array[23184] <= 3'b111;
      // memory_array[23185] <= 3'b110;
      // memory_array[23186] <= 3'b110;
      // memory_array[23187] <= 3'b110;
      // memory_array[23188] <= 3'b000;
      // memory_array[23189] <= 3'b000;
      // memory_array[23190] <= 3'b000;
      // memory_array[23191] <= 3'b101;
      // memory_array[23192] <= 3'b101;
      // memory_array[23193] <= 3'b101;
      // memory_array[23194] <= 3'b000;
      // memory_array[23195] <= 3'b101;
      // memory_array[23196] <= 3'b101;
      // memory_array[23197] <= 3'b110;
      // memory_array[23198] <= 3'b101;
      // memory_array[23199] <= 3'b101;
      // memory_array[23200] <= 3'b101;
      // memory_array[23201] <= 3'b110;
      // memory_array[23202] <= 3'b110;
      // memory_array[23203] <= 3'b000;
      // memory_array[23204] <= 3'b000;
      // memory_array[23205] <= 3'b110;
      // memory_array[23206] <= 3'b110;
      // memory_array[23207] <= 3'b101;
      // memory_array[23208] <= 3'b101;
      // memory_array[23209] <= 3'b000;
      // memory_array[23210] <= 3'b000;
      // memory_array[23211] <= 3'b110;
      // memory_array[23212] <= 3'b110;
      // memory_array[23213] <= 3'b110;
      // memory_array[23214] <= 3'b110;
      // memory_array[23215] <= 3'b110;
      // memory_array[23216] <= 3'b110;
      // memory_array[23217] <= 3'b110;
      // memory_array[23218] <= 3'b111;
      // memory_array[23219] <= 3'b111;
      // memory_array[23220] <= 3'b110;
      // memory_array[23221] <= 3'b000;
      // memory_array[23222] <= 3'b110;
      // memory_array[23223] <= 3'b000;
      // memory_array[23224] <= 3'b111;
      // memory_array[23225] <= 3'b111;
      // memory_array[23226] <= 3'b111;
      // memory_array[23227] <= 3'b000;
      // memory_array[23228] <= 3'b111;
      // memory_array[23229] <= 3'b111;
      // memory_array[23230] <= 3'b110;
      // memory_array[23231] <= 3'b110;
      // memory_array[23232] <= 3'b000;
      // memory_array[23233] <= 3'b111;
      // memory_array[23234] <= 3'b110;
      // memory_array[23235] <= 3'b110;
      // memory_array[23236] <= 3'b110;
      // memory_array[23237] <= 3'b111;
      // memory_array[23238] <= 3'b111;
      // memory_array[23239] <= 3'b111;
      // memory_array[23240] <= 3'b111;
      // memory_array[23241] <= 3'b000;
      // memory_array[23242] <= 3'b110;
      // memory_array[23243] <= 3'b000;
      // memory_array[23244] <= 3'b111;
      // memory_array[23245] <= 3'b000;
      // memory_array[23246] <= 3'b111;
      // memory_array[23247] <= 3'b000;
      // memory_array[23248] <= 3'b000;
      // memory_array[23249] <= 3'b101;
      // memory_array[23250] <= 3'b000;
      // memory_array[23251] <= 3'b000;
      // memory_array[23252] <= 3'b000;
      // memory_array[23253] <= 3'b000;
      // memory_array[23254] <= 3'b000;
      // memory_array[23255] <= 3'b101;
      // memory_array[23256] <= 3'b101;
      // memory_array[23257] <= 3'b101;
      // memory_array[23258] <= 3'b000;
      // memory_array[23259] <= 3'b000;
      // memory_array[23260] <= 3'b000;
      // memory_array[23261] <= 3'b000;
      // memory_array[23262] <= 3'b000;
      // memory_array[23263] <= 3'b000;
      // memory_array[23264] <= 3'b000;
      // memory_array[23265] <= 3'b000;
      // memory_array[23266] <= 3'b000;
      // memory_array[23267] <= 3'b000;
      // memory_array[23268] <= 3'b000;
      // memory_array[23269] <= 3'b000;
      // memory_array[23270] <= 3'b000;
      // memory_array[23271] <= 3'b000;
      // memory_array[23272] <= 3'b000;
      // memory_array[23273] <= 3'b000;
      // memory_array[23274] <= 3'b000;
      // memory_array[23275] <= 3'b000;
      // memory_array[23276] <= 3'b000;
      // memory_array[23277] <= 3'b000;
      // memory_array[23278] <= 3'b000;
      // memory_array[23279] <= 3'b000;
      // memory_array[23280] <= 3'b101;
      // memory_array[23281] <= 3'b000;
      // memory_array[23282] <= 3'b000;
      // memory_array[23283] <= 3'b000;
      // memory_array[23284] <= 3'b000;
      // memory_array[23285] <= 3'b000;
      // memory_array[23286] <= 3'b000;
      // memory_array[23287] <= 3'b000;
      // memory_array[23288] <= 3'b000;
      // memory_array[23289] <= 3'b000;
      // memory_array[23290] <= 3'b101;
      // memory_array[23291] <= 3'b101;
      // memory_array[23292] <= 3'b101;
      // memory_array[23293] <= 3'b000;
      // memory_array[23294] <= 3'b000;
      // memory_array[23295] <= 3'b000;
      // memory_array[23296] <= 3'b000;
      // memory_array[23297] <= 3'b000;
      // memory_array[23298] <= 3'b000;
      // memory_array[23299] <= 3'b000;
      // memory_array[23300] <= 3'b000;
      // memory_array[23301] <= 3'b000;
      // memory_array[23302] <= 3'b000;
      // memory_array[23303] <= 3'b000;
      // memory_array[23304] <= 3'b000;
      // memory_array[23305] <= 3'b000;
      // memory_array[23306] <= 3'b000;
      // memory_array[23307] <= 3'b101;
      // memory_array[23308] <= 3'b101;
      // memory_array[23309] <= 3'b101;
      // memory_array[23310] <= 3'b000;
      // memory_array[23311] <= 3'b101;
      // memory_array[23312] <= 3'b101;
      // memory_array[23313] <= 3'b101;
      // memory_array[23314] <= 3'b101;
      // memory_array[23315] <= 3'b101;
      // memory_array[23316] <= 3'b101;
      // memory_array[23317] <= 3'b101;
      // memory_array[23318] <= 3'b000;
      // memory_array[23319] <= 3'b000;
      // memory_array[23320] <= 3'b000;
      // memory_array[23321] <= 3'b000;
      // memory_array[23322] <= 3'b000;
      // memory_array[23323] <= 3'b000;
      // memory_array[23324] <= 3'b000;
      // memory_array[23325] <= 3'b000;
      // memory_array[23326] <= 3'b000;
      // memory_array[23327] <= 3'b000;
      // memory_array[23328] <= 3'b000;
      // memory_array[23329] <= 3'b000;
      // memory_array[23330] <= 3'b000;
      // memory_array[23331] <= 3'b000;
      // memory_array[23332] <= 3'b000;
      // memory_array[23333] <= 3'b000;
      // memory_array[23334] <= 3'b000;
      // memory_array[23335] <= 3'b000;
      // memory_array[23336] <= 3'b101;
      // memory_array[23337] <= 3'b000;
      // memory_array[23338] <= 3'b000;
      // memory_array[23339] <= 3'b000;
      // memory_array[23340] <= 3'b000;
      // memory_array[23341] <= 3'b000;
      // memory_array[23342] <= 3'b000;
      // memory_array[23343] <= 3'b000;
      // memory_array[23344] <= 3'b000;
      // memory_array[23345] <= 3'b101;
      // memory_array[23346] <= 3'b000;
      // memory_array[23347] <= 3'b000;
      // memory_array[23348] <= 3'b000;
      // memory_array[23349] <= 3'b000;
      // memory_array[23350] <= 3'b111;
      // memory_array[23351] <= 3'b111;
      // memory_array[23352] <= 3'b000;
      // memory_array[23353] <= 3'b111;
      // memory_array[23354] <= 3'b111;
      // memory_array[23355] <= 3'b101;
      // memory_array[23356] <= 3'b110;
      // memory_array[23357] <= 3'b110;
      // memory_array[23358] <= 3'b110;
      // memory_array[23359] <= 3'b110;
      // memory_array[23360] <= 3'b110;
      // memory_array[23361] <= 3'b111;
      // memory_array[23362] <= 3'b111;
      // memory_array[23363] <= 3'b111;
      // memory_array[23364] <= 3'b111;
      // memory_array[23365] <= 3'b111;
      // memory_array[23366] <= 3'b110;
      // memory_array[23367] <= 3'b111;
      // memory_array[23368] <= 3'b111;
      // memory_array[23369] <= 3'b111;
      // memory_array[23370] <= 3'b111;
      // memory_array[23371] <= 3'b111;
      // memory_array[23372] <= 3'b000;
      // memory_array[23373] <= 3'b110;
      // memory_array[23374] <= 3'b000;
      // memory_array[23375] <= 3'b111;
      // memory_array[23376] <= 3'b111;
      // memory_array[23377] <= 3'b111;
      // memory_array[23378] <= 3'b111;
      // memory_array[23379] <= 3'b110;
      // memory_array[23380] <= 3'b110;
      // memory_array[23381] <= 3'b110;
      // memory_array[23382] <= 3'b110;
      // memory_array[23383] <= 3'b111;
      // memory_array[23384] <= 3'b111;
      // memory_array[23385] <= 3'b110;
      // memory_array[23386] <= 3'b110;
      // memory_array[23387] <= 3'b110;
      // memory_array[23388] <= 3'b111;
      // memory_array[23389] <= 3'b000;
      // memory_array[23390] <= 3'b000;
      // memory_array[23391] <= 3'b101;
      // memory_array[23392] <= 3'b110;
      // memory_array[23393] <= 3'b000;
      // memory_array[23394] <= 3'b000;
      // memory_array[23395] <= 3'b110;
      // memory_array[23396] <= 3'b110;
      // memory_array[23397] <= 3'b110;
      // memory_array[23398] <= 3'b000;
      // memory_array[23399] <= 3'b101;
      // memory_array[23400] <= 3'b000;
      // memory_array[23401] <= 3'b000;
      // memory_array[23402] <= 3'b000;
      // memory_array[23403] <= 3'b110;
      // memory_array[23404] <= 3'b110;
      // memory_array[23405] <= 3'b000;
      // memory_array[23406] <= 3'b000;
      // memory_array[23407] <= 3'b000;
      // memory_array[23408] <= 3'b101;
      // memory_array[23409] <= 3'b000;
      // memory_array[23410] <= 3'b000;
      // memory_array[23411] <= 3'b110;
      // memory_array[23412] <= 3'b111;
      // memory_array[23413] <= 3'b110;
      // memory_array[23414] <= 3'b110;
      // memory_array[23415] <= 3'b110;
      // memory_array[23416] <= 3'b111;
      // memory_array[23417] <= 3'b110;
      // memory_array[23418] <= 3'b110;
      // memory_array[23419] <= 3'b110;
      // memory_array[23420] <= 3'b110;
      // memory_array[23421] <= 3'b000;
      // memory_array[23422] <= 3'b000;
      // memory_array[23423] <= 3'b000;
      // memory_array[23424] <= 3'b111;
      // memory_array[23425] <= 3'b111;
      // memory_array[23426] <= 3'b111;
      // memory_array[23427] <= 3'b000;
      // memory_array[23428] <= 3'b110;
      // memory_array[23429] <= 3'b110;
      // memory_array[23430] <= 3'b110;
      // memory_array[23431] <= 3'b110;
      // memory_array[23432] <= 3'b000;
      // memory_array[23433] <= 3'b110;
      // memory_array[23434] <= 3'b110;
      // memory_array[23435] <= 3'b111;
      // memory_array[23436] <= 3'b111;
      // memory_array[23437] <= 3'b111;
      // memory_array[23438] <= 3'b111;
      // memory_array[23439] <= 3'b111;
      // memory_array[23440] <= 3'b111;
      // memory_array[23441] <= 3'b111;
      // memory_array[23442] <= 3'b000;
      // memory_array[23443] <= 3'b000;
      // memory_array[23444] <= 3'b111;
      // memory_array[23445] <= 3'b111;
      // memory_array[23446] <= 3'b000;
      // memory_array[23447] <= 3'b111;
      // memory_array[23448] <= 3'b111;
      // memory_array[23449] <= 3'b101;
      // memory_array[23450] <= 3'b000;
      // memory_array[23451] <= 3'b000;
      // memory_array[23452] <= 3'b000;
      // memory_array[23453] <= 3'b101;
      // memory_array[23454] <= 3'b101;
      // memory_array[23455] <= 3'b000;
      // memory_array[23456] <= 3'b000;
      // memory_array[23457] <= 3'b000;
      // memory_array[23458] <= 3'b101;
      // memory_array[23459] <= 3'b000;
      // memory_array[23460] <= 3'b000;
      // memory_array[23461] <= 3'b000;
      // memory_array[23462] <= 3'b000;
      // memory_array[23463] <= 3'b000;
      // memory_array[23464] <= 3'b000;
      // memory_array[23465] <= 3'b000;
      // memory_array[23466] <= 3'b000;
      // memory_array[23467] <= 3'b000;
      // memory_array[23468] <= 3'b000;
      // memory_array[23469] <= 3'b000;
      // memory_array[23470] <= 3'b000;
      // memory_array[23471] <= 3'b000;
      // memory_array[23472] <= 3'b000;
      // memory_array[23473] <= 3'b101;
      // memory_array[23474] <= 3'b101;
      // memory_array[23475] <= 3'b000;
      // memory_array[23476] <= 3'b000;
      // memory_array[23477] <= 3'b000;
      // memory_array[23478] <= 3'b000;
      // memory_array[23479] <= 3'b000;
      // memory_array[23480] <= 3'b000;
      // memory_array[23481] <= 3'b000;
      // memory_array[23482] <= 3'b000;
      // memory_array[23483] <= 3'b000;
      // memory_array[23484] <= 3'b000;
      // memory_array[23485] <= 3'b000;
      // memory_array[23486] <= 3'b000;
      // memory_array[23487] <= 3'b000;
      // memory_array[23488] <= 3'b000;
      // memory_array[23489] <= 3'b101;
      // memory_array[23490] <= 3'b000;
      // memory_array[23491] <= 3'b000;
      // memory_array[23492] <= 3'b000;
      // memory_array[23493] <= 3'b101;
      // memory_array[23494] <= 3'b000;
      // memory_array[23495] <= 3'b000;
      // memory_array[23496] <= 3'b000;
      // memory_array[23497] <= 3'b000;
      // memory_array[23498] <= 3'b101;
      // memory_array[23499] <= 3'b000;
      // memory_array[23500] <= 3'b000;
      // memory_array[23501] <= 3'b000;
      // memory_array[23502] <= 3'b101;
      // memory_array[23503] <= 3'b101;
      // memory_array[23504] <= 3'b101;
      // memory_array[23505] <= 3'b101;
      // memory_array[23506] <= 3'b101;
      // memory_array[23507] <= 3'b101;
      // memory_array[23508] <= 3'b101;
      // memory_array[23509] <= 3'b101;
      // memory_array[23510] <= 3'b101;
      // memory_array[23511] <= 3'b101;
      // memory_array[23512] <= 3'b101;
      // memory_array[23513] <= 3'b101;
      // memory_array[23514] <= 3'b101;
      // memory_array[23515] <= 3'b101;
      // memory_array[23516] <= 3'b101;
      // memory_array[23517] <= 3'b101;
      // memory_array[23518] <= 3'b101;
      // memory_array[23519] <= 3'b101;
      // memory_array[23520] <= 3'b000;
      // memory_array[23521] <= 3'b000;
      // memory_array[23522] <= 3'b000;
      // memory_array[23523] <= 3'b101;
      // memory_array[23524] <= 3'b000;
      // memory_array[23525] <= 3'b000;
      // memory_array[23526] <= 3'b000;
      // memory_array[23527] <= 3'b000;
      // memory_array[23528] <= 3'b000;
      // memory_array[23529] <= 3'b000;
      // memory_array[23530] <= 3'b000;
      // memory_array[23531] <= 3'b000;
      // memory_array[23532] <= 3'b000;
      // memory_array[23533] <= 3'b000;
      // memory_array[23534] <= 3'b000;
      // memory_array[23535] <= 3'b000;
      // memory_array[23536] <= 3'b000;
      // memory_array[23537] <= 3'b000;
      // memory_array[23538] <= 3'b101;
      // memory_array[23539] <= 3'b101;
      // memory_array[23540] <= 3'b000;
      // memory_array[23541] <= 3'b000;
      // memory_array[23542] <= 3'b000;
      // memory_array[23543] <= 3'b000;
      // memory_array[23544] <= 3'b000;
      // memory_array[23545] <= 3'b000;
      // memory_array[23546] <= 3'b000;
      // memory_array[23547] <= 3'b000;
      // memory_array[23548] <= 3'b000;
      // memory_array[23549] <= 3'b000;
      // memory_array[23550] <= 3'b111;
      // memory_array[23551] <= 3'b111;
      // memory_array[23552] <= 3'b111;
      // memory_array[23553] <= 3'b111;
      // memory_array[23554] <= 3'b111;
      // memory_array[23555] <= 3'b101;
      // memory_array[23556] <= 3'b110;
      // memory_array[23557] <= 3'b000;
      // memory_array[23558] <= 3'b110;
      // memory_array[23559] <= 3'b000;
      // memory_array[23560] <= 3'b000;
      // memory_array[23561] <= 3'b111;
      // memory_array[23562] <= 3'b111;
      // memory_array[23563] <= 3'b111;
      // memory_array[23564] <= 3'b111;
      // memory_array[23565] <= 3'b111;
      // memory_array[23566] <= 3'b110;
      // memory_array[23567] <= 3'b000;
      // memory_array[23568] <= 3'b111;
      // memory_array[23569] <= 3'b111;
      // memory_array[23570] <= 3'b111;
      // memory_array[23571] <= 3'b111;
      // memory_array[23572] <= 3'b111;
      // memory_array[23573] <= 3'b000;
      // memory_array[23574] <= 3'b000;
      // memory_array[23575] <= 3'b111;
      // memory_array[23576] <= 3'b111;
      // memory_array[23577] <= 3'b111;
      // memory_array[23578] <= 3'b111;
      // memory_array[23579] <= 3'b110;
      // memory_array[23580] <= 3'b111;
      // memory_array[23581] <= 3'b111;
      // memory_array[23582] <= 3'b111;
      // memory_array[23583] <= 3'b110;
      // memory_array[23584] <= 3'b110;
      // memory_array[23585] <= 3'b111;
      // memory_array[23586] <= 3'b111;
      // memory_array[23587] <= 3'b111;
      // memory_array[23588] <= 3'b110;
      // memory_array[23589] <= 3'b000;
      // memory_array[23590] <= 3'b000;
      // memory_array[23591] <= 3'b101;
      // memory_array[23592] <= 3'b000;
      // memory_array[23593] <= 3'b110;
      // memory_array[23594] <= 3'b110;
      // memory_array[23595] <= 3'b000;
      // memory_array[23596] <= 3'b000;
      // memory_array[23597] <= 3'b000;
      // memory_array[23598] <= 3'b110;
      // memory_array[23599] <= 3'b110;
      // memory_array[23600] <= 3'b101;
      // memory_array[23601] <= 3'b101;
      // memory_array[23602] <= 3'b101;
      // memory_array[23603] <= 3'b101;
      // memory_array[23604] <= 3'b101;
      // memory_array[23605] <= 3'b101;
      // memory_array[23606] <= 3'b101;
      // memory_array[23607] <= 3'b101;
      // memory_array[23608] <= 3'b101;
      // memory_array[23609] <= 3'b000;
      // memory_array[23610] <= 3'b000;
      // memory_array[23611] <= 3'b110;
      // memory_array[23612] <= 3'b110;
      // memory_array[23613] <= 3'b111;
      // memory_array[23614] <= 3'b111;
      // memory_array[23615] <= 3'b110;
      // memory_array[23616] <= 3'b110;
      // memory_array[23617] <= 3'b110;
      // memory_array[23618] <= 3'b110;
      // memory_array[23619] <= 3'b110;
      // memory_array[23620] <= 3'b110;
      // memory_array[23621] <= 3'b000;
      // memory_array[23622] <= 3'b110;
      // memory_array[23623] <= 3'b000;
      // memory_array[23624] <= 3'b111;
      // memory_array[23625] <= 3'b111;
      // memory_array[23626] <= 3'b111;
      // memory_array[23627] <= 3'b000;
      // memory_array[23628] <= 3'b110;
      // memory_array[23629] <= 3'b110;
      // memory_array[23630] <= 3'b110;
      // memory_array[23631] <= 3'b110;
      // memory_array[23632] <= 3'b000;
      // memory_array[23633] <= 3'b110;
      // memory_array[23634] <= 3'b111;
      // memory_array[23635] <= 3'b110;
      // memory_array[23636] <= 3'b000;
      // memory_array[23637] <= 3'b111;
      // memory_array[23638] <= 3'b111;
      // memory_array[23639] <= 3'b111;
      // memory_array[23640] <= 3'b111;
      // memory_array[23641] <= 3'b111;
      // memory_array[23642] <= 3'b111;
      // memory_array[23643] <= 3'b111;
      // memory_array[23644] <= 3'b111;
      // memory_array[23645] <= 3'b111;
      // memory_array[23646] <= 3'b111;
      // memory_array[23647] <= 3'b111;
      // memory_array[23648] <= 3'b111;
      // memory_array[23649] <= 3'b101;
      // memory_array[23650] <= 3'b000;
      // memory_array[23651] <= 3'b110;
      // memory_array[23652] <= 3'b101;
      // memory_array[23653] <= 3'b000;
      // memory_array[23654] <= 3'b000;
      // memory_array[23655] <= 3'b000;
      // memory_array[23656] <= 3'b101;
      // memory_array[23657] <= 3'b101;
      // memory_array[23658] <= 3'b000;
      // memory_array[23659] <= 3'b000;
      // memory_array[23660] <= 3'b000;
      // memory_array[23661] <= 3'b000;
      // memory_array[23662] <= 3'b000;
      // memory_array[23663] <= 3'b000;
      // memory_array[23664] <= 3'b000;
      // memory_array[23665] <= 3'b000;
      // memory_array[23666] <= 3'b000;
      // memory_array[23667] <= 3'b000;
      // memory_array[23668] <= 3'b000;
      // memory_array[23669] <= 3'b000;
      // memory_array[23670] <= 3'b101;
      // memory_array[23671] <= 3'b101;
      // memory_array[23672] <= 3'b101;
      // memory_array[23673] <= 3'b000;
      // memory_array[23674] <= 3'b000;
      // memory_array[23675] <= 3'b000;
      // memory_array[23676] <= 3'b101;
      // memory_array[23677] <= 3'b101;
      // memory_array[23678] <= 3'b000;
      // memory_array[23679] <= 3'b000;
      // memory_array[23680] <= 3'b000;
      // memory_array[23681] <= 3'b000;
      // memory_array[23682] <= 3'b101;
      // memory_array[23683] <= 3'b000;
      // memory_array[23684] <= 3'b000;
      // memory_array[23685] <= 3'b000;
      // memory_array[23686] <= 3'b000;
      // memory_array[23687] <= 3'b000;
      // memory_array[23688] <= 3'b000;
      // memory_array[23689] <= 3'b000;
      // memory_array[23690] <= 3'b101;
      // memory_array[23691] <= 3'b101;
      // memory_array[23692] <= 3'b101;
      // memory_array[23693] <= 3'b000;
      // memory_array[23694] <= 3'b000;
      // memory_array[23695] <= 3'b000;
      // memory_array[23696] <= 3'b000;
      // memory_array[23697] <= 3'b101;
      // memory_array[23698] <= 3'b000;
      // memory_array[23699] <= 3'b000;
      // memory_array[23700] <= 3'b000;
      // memory_array[23701] <= 3'b101;
      // memory_array[23702] <= 3'b101;
      // memory_array[23703] <= 3'b101;
      // memory_array[23704] <= 3'b101;
      // memory_array[23705] <= 3'b101;
      // memory_array[23706] <= 3'b101;
      // memory_array[23707] <= 3'b101;
      // memory_array[23708] <= 3'b101;
      // memory_array[23709] <= 3'b101;
      // memory_array[23710] <= 3'b101;
      // memory_array[23711] <= 3'b101;
      // memory_array[23712] <= 3'b101;
      // memory_array[23713] <= 3'b000;
      // memory_array[23714] <= 3'b000;
      // memory_array[23715] <= 3'b101;
      // memory_array[23716] <= 3'b000;
      // memory_array[23717] <= 3'b000;
      // memory_array[23718] <= 3'b000;
      // memory_array[23719] <= 3'b000;
      // memory_array[23720] <= 3'b101;
      // memory_array[23721] <= 3'b000;
      // memory_array[23722] <= 3'b000;
      // memory_array[23723] <= 3'b000;
      // memory_array[23724] <= 3'b000;
      // memory_array[23725] <= 3'b101;
      // memory_array[23726] <= 3'b000;
      // memory_array[23727] <= 3'b000;
      // memory_array[23728] <= 3'b000;
      // memory_array[23729] <= 3'b000;
      // memory_array[23730] <= 3'b000;
      // memory_array[23731] <= 3'b000;
      // memory_array[23732] <= 3'b000;
      // memory_array[23733] <= 3'b000;
      // memory_array[23734] <= 3'b000;
      // memory_array[23735] <= 3'b000;
      // memory_array[23736] <= 3'b000;
      // memory_array[23737] <= 3'b101;
      // memory_array[23738] <= 3'b000;
      // memory_array[23739] <= 3'b000;
      // memory_array[23740] <= 3'b000;
      // memory_array[23741] <= 3'b101;
      // memory_array[23742] <= 3'b101;
      // memory_array[23743] <= 3'b000;
      // memory_array[23744] <= 3'b000;
      // memory_array[23745] <= 3'b000;
      // memory_array[23746] <= 3'b101;
      // memory_array[23747] <= 3'b000;
      // memory_array[23748] <= 3'b000;
      // memory_array[23749] <= 3'b000;
      // memory_array[23750] <= 3'b111;
      // memory_array[23751] <= 3'b111;
      // memory_array[23752] <= 3'b111;
      // memory_array[23753] <= 3'b111;
      // memory_array[23754] <= 3'b111;
      // memory_array[23755] <= 3'b101;
      // memory_array[23756] <= 3'b110;
      // memory_array[23757] <= 3'b110;
      // memory_array[23758] <= 3'b000;
      // memory_array[23759] <= 3'b111;
      // memory_array[23760] <= 3'b111;
      // memory_array[23761] <= 3'b111;
      // memory_array[23762] <= 3'b111;
      // memory_array[23763] <= 3'b111;
      // memory_array[23764] <= 3'b111;
      // memory_array[23765] <= 3'b111;
      // memory_array[23766] <= 3'b110;
      // memory_array[23767] <= 3'b000;
      // memory_array[23768] <= 3'b111;
      // memory_array[23769] <= 3'b111;
      // memory_array[23770] <= 3'b111;
      // memory_array[23771] <= 3'b111;
      // memory_array[23772] <= 3'b111;
      // memory_array[23773] <= 3'b111;
      // memory_array[23774] <= 3'b000;
      // memory_array[23775] <= 3'b111;
      // memory_array[23776] <= 3'b111;
      // memory_array[23777] <= 3'b111;
      // memory_array[23778] <= 3'b111;
      // memory_array[23779] <= 3'b111;
      // memory_array[23780] <= 3'b110;
      // memory_array[23781] <= 3'b110;
      // memory_array[23782] <= 3'b110;
      // memory_array[23783] <= 3'b110;
      // memory_array[23784] <= 3'b110;
      // memory_array[23785] <= 3'b110;
      // memory_array[23786] <= 3'b110;
      // memory_array[23787] <= 3'b110;
      // memory_array[23788] <= 3'b110;
      // memory_array[23789] <= 3'b000;
      // memory_array[23790] <= 3'b000;
      // memory_array[23791] <= 3'b101;
      // memory_array[23792] <= 3'b101;
      // memory_array[23793] <= 3'b101;
      // memory_array[23794] <= 3'b101;
      // memory_array[23795] <= 3'b101;
      // memory_array[23796] <= 3'b101;
      // memory_array[23797] <= 3'b101;
      // memory_array[23798] <= 3'b101;
      // memory_array[23799] <= 3'b101;
      // memory_array[23800] <= 3'b101;
      // memory_array[23801] <= 3'b101;
      // memory_array[23802] <= 3'b101;
      // memory_array[23803] <= 3'b101;
      // memory_array[23804] <= 3'b101;
      // memory_array[23805] <= 3'b101;
      // memory_array[23806] <= 3'b101;
      // memory_array[23807] <= 3'b101;
      // memory_array[23808] <= 3'b101;
      // memory_array[23809] <= 3'b000;
      // memory_array[23810] <= 3'b000;
      // memory_array[23811] <= 3'b110;
      // memory_array[23812] <= 3'b110;
      // memory_array[23813] <= 3'b111;
      // memory_array[23814] <= 3'b111;
      // memory_array[23815] <= 3'b110;
      // memory_array[23816] <= 3'b110;
      // memory_array[23817] <= 3'b110;
      // memory_array[23818] <= 3'b110;
      // memory_array[23819] <= 3'b110;
      // memory_array[23820] <= 3'b110;
      // memory_array[23821] <= 3'b000;
      // memory_array[23822] <= 3'b110;
      // memory_array[23823] <= 3'b000;
      // memory_array[23824] <= 3'b111;
      // memory_array[23825] <= 3'b111;
      // memory_array[23826] <= 3'b111;
      // memory_array[23827] <= 3'b000;
      // memory_array[23828] <= 3'b110;
      // memory_array[23829] <= 3'b110;
      // memory_array[23830] <= 3'b110;
      // memory_array[23831] <= 3'b110;
      // memory_array[23832] <= 3'b000;
      // memory_array[23833] <= 3'b110;
      // memory_array[23834] <= 3'b111;
      // memory_array[23835] <= 3'b110;
      // memory_array[23836] <= 3'b111;
      // memory_array[23837] <= 3'b111;
      // memory_array[23838] <= 3'b111;
      // memory_array[23839] <= 3'b111;
      // memory_array[23840] <= 3'b000;
      // memory_array[23841] <= 3'b000;
      // memory_array[23842] <= 3'b110;
      // memory_array[23843] <= 3'b000;
      // memory_array[23844] <= 3'b111;
      // memory_array[23845] <= 3'b111;
      // memory_array[23846] <= 3'b111;
      // memory_array[23847] <= 3'b111;
      // memory_array[23848] <= 3'b111;
      // memory_array[23849] <= 3'b101;
      // memory_array[23850] <= 3'b000;
      // memory_array[23851] <= 3'b000;
      // memory_array[23852] <= 3'b000;
      // memory_array[23853] <= 3'b000;
      // memory_array[23854] <= 3'b000;
      // memory_array[23855] <= 3'b101;
      // memory_array[23856] <= 3'b000;
      // memory_array[23857] <= 3'b000;
      // memory_array[23858] <= 3'b000;
      // memory_array[23859] <= 3'b000;
      // memory_array[23860] <= 3'b000;
      // memory_array[23861] <= 3'b000;
      // memory_array[23862] <= 3'b000;
      // memory_array[23863] <= 3'b000;
      // memory_array[23864] <= 3'b000;
      // memory_array[23865] <= 3'b000;
      // memory_array[23866] <= 3'b000;
      // memory_array[23867] <= 3'b101;
      // memory_array[23868] <= 3'b000;
      // memory_array[23869] <= 3'b000;
      // memory_array[23870] <= 3'b101;
      // memory_array[23871] <= 3'b101;
      // memory_array[23872] <= 3'b000;
      // memory_array[23873] <= 3'b000;
      // memory_array[23874] <= 3'b000;
      // memory_array[23875] <= 3'b000;
      // memory_array[23876] <= 3'b000;
      // memory_array[23877] <= 3'b101;
      // memory_array[23878] <= 3'b000;
      // memory_array[23879] <= 3'b000;
      // memory_array[23880] <= 3'b000;
      // memory_array[23881] <= 3'b000;
      // memory_array[23882] <= 3'b000;
      // memory_array[23883] <= 3'b000;
      // memory_array[23884] <= 3'b000;
      // memory_array[23885] <= 3'b000;
      // memory_array[23886] <= 3'b101;
      // memory_array[23887] <= 3'b000;
      // memory_array[23888] <= 3'b000;
      // memory_array[23889] <= 3'b000;
      // memory_array[23890] <= 3'b000;
      // memory_array[23891] <= 3'b000;
      // memory_array[23892] <= 3'b000;
      // memory_array[23893] <= 3'b000;
      // memory_array[23894] <= 3'b000;
      // memory_array[23895] <= 3'b000;
      // memory_array[23896] <= 3'b000;
      // memory_array[23897] <= 3'b000;
      // memory_array[23898] <= 3'b000;
      // memory_array[23899] <= 3'b000;
      // memory_array[23900] <= 3'b000;
      // memory_array[23901] <= 3'b000;
      // memory_array[23902] <= 3'b000;
      // memory_array[23903] <= 3'b000;
      // memory_array[23904] <= 3'b000;
      // memory_array[23905] <= 3'b000;
      // memory_array[23906] <= 3'b000;
      // memory_array[23907] <= 3'b000;
      // memory_array[23908] <= 3'b000;
      // memory_array[23909] <= 3'b101;
      // memory_array[23910] <= 3'b000;
      // memory_array[23911] <= 3'b101;
      // memory_array[23912] <= 3'b000;
      // memory_array[23913] <= 3'b000;
      // memory_array[23914] <= 3'b000;
      // memory_array[23915] <= 3'b101;
      // memory_array[23916] <= 3'b000;
      // memory_array[23917] <= 3'b101;
      // memory_array[23918] <= 3'b000;
      // memory_array[23919] <= 3'b000;
      // memory_array[23920] <= 3'b000;
      // memory_array[23921] <= 3'b000;
      // memory_array[23922] <= 3'b000;
      // memory_array[23923] <= 3'b000;
      // memory_array[23924] <= 3'b000;
      // memory_array[23925] <= 3'b000;
      // memory_array[23926] <= 3'b000;
      // memory_array[23927] <= 3'b000;
      // memory_array[23928] <= 3'b000;
      // memory_array[23929] <= 3'b000;
      // memory_array[23930] <= 3'b000;
      // memory_array[23931] <= 3'b000;
      // memory_array[23932] <= 3'b000;
      // memory_array[23933] <= 3'b000;
      // memory_array[23934] <= 3'b000;
      // memory_array[23935] <= 3'b000;
      // memory_array[23936] <= 3'b101;
      // memory_array[23937] <= 3'b101;
      // memory_array[23938] <= 3'b000;
      // memory_array[23939] <= 3'b000;
      // memory_array[23940] <= 3'b000;
      // memory_array[23941] <= 3'b101;
      // memory_array[23942] <= 3'b101;
      // memory_array[23943] <= 3'b000;
      // memory_array[23944] <= 3'b000;
      // memory_array[23945] <= 3'b101;
      // memory_array[23946] <= 3'b000;
      // memory_array[23947] <= 3'b000;
      // memory_array[23948] <= 3'b000;
      // memory_array[23949] <= 3'b000;
      // memory_array[23950] <= 3'b111;
      // memory_array[23951] <= 3'b111;
      // memory_array[23952] <= 3'b111;
      // memory_array[23953] <= 3'b111;
      // memory_array[23954] <= 3'b111;
      // memory_array[23955] <= 3'b101;
      // memory_array[23956] <= 3'b110;
      // memory_array[23957] <= 3'b110;
      // memory_array[23958] <= 3'b000;
      // memory_array[23959] <= 3'b000;
      // memory_array[23960] <= 3'b000;
      // memory_array[23961] <= 3'b000;
      // memory_array[23962] <= 3'b111;
      // memory_array[23963] <= 3'b111;
      // memory_array[23964] <= 3'b111;
      // memory_array[23965] <= 3'b111;
      // memory_array[23966] <= 3'b000;
      // memory_array[23967] <= 3'b110;
      // memory_array[23968] <= 3'b000;
      // memory_array[23969] <= 3'b111;
      // memory_array[23970] <= 3'b111;
      // memory_array[23971] <= 3'b111;
      // memory_array[23972] <= 3'b111;
      // memory_array[23973] <= 3'b111;
      // memory_array[23974] <= 3'b111;
      // memory_array[23975] <= 3'b111;
      // memory_array[23976] <= 3'b111;
      // memory_array[23977] <= 3'b111;
      // memory_array[23978] <= 3'b111;
      // memory_array[23979] <= 3'b111;
      // memory_array[23980] <= 3'b110;
      // memory_array[23981] <= 3'b110;
      // memory_array[23982] <= 3'b110;
      // memory_array[23983] <= 3'b110;
      // memory_array[23984] <= 3'b110;
      // memory_array[23985] <= 3'b110;
      // memory_array[23986] <= 3'b110;
      // memory_array[23987] <= 3'b110;
      // memory_array[23988] <= 3'b110;
      // memory_array[23989] <= 3'b000;
      // memory_array[23990] <= 3'b000;
      // memory_array[23991] <= 3'b101;
      // memory_array[23992] <= 3'b101;
      // memory_array[23993] <= 3'b101;
      // memory_array[23994] <= 3'b101;
      // memory_array[23995] <= 3'b101;
      // memory_array[23996] <= 3'b101;
      // memory_array[23997] <= 3'b101;
      // memory_array[23998] <= 3'b101;
      // memory_array[23999] <= 3'b101;
      // memory_array[24000] <= 3'b000;
      // memory_array[24001] <= 3'b000;
      // memory_array[24002] <= 3'b000;
      // memory_array[24003] <= 3'b110;
      // memory_array[24004] <= 3'b110;
      // memory_array[24005] <= 3'b000;
      // memory_array[24006] <= 3'b000;
      // memory_array[24007] <= 3'b000;
      // memory_array[24008] <= 3'b101;
      // memory_array[24009] <= 3'b000;
      // memory_array[24010] <= 3'b000;
      // memory_array[24011] <= 3'b110;
      // memory_array[24012] <= 3'b111;
      // memory_array[24013] <= 3'b110;
      // memory_array[24014] <= 3'b110;
      // memory_array[24015] <= 3'b110;
      // memory_array[24016] <= 3'b111;
      // memory_array[24017] <= 3'b110;
      // memory_array[24018] <= 3'b110;
      // memory_array[24019] <= 3'b110;
      // memory_array[24020] <= 3'b110;
      // memory_array[24021] <= 3'b000;
      // memory_array[24022] <= 3'b000;
      // memory_array[24023] <= 3'b000;
      // memory_array[24024] <= 3'b111;
      // memory_array[24025] <= 3'b111;
      // memory_array[24026] <= 3'b111;
      // memory_array[24027] <= 3'b000;
      // memory_array[24028] <= 3'b110;
      // memory_array[24029] <= 3'b110;
      // memory_array[24030] <= 3'b110;
      // memory_array[24031] <= 3'b110;
      // memory_array[24032] <= 3'b000;
      // memory_array[24033] <= 3'b110;
      // memory_array[24034] <= 3'b000;
      // memory_array[24035] <= 3'b000;
      // memory_array[24036] <= 3'b111;
      // memory_array[24037] <= 3'b000;
      // memory_array[24038] <= 3'b000;
      // memory_array[24039] <= 3'b000;
      // memory_array[24040] <= 3'b000;
      // memory_array[24041] <= 3'b000;
      // memory_array[24042] <= 3'b000;
      // memory_array[24043] <= 3'b110;
      // memory_array[24044] <= 3'b111;
      // memory_array[24045] <= 3'b111;
      // memory_array[24046] <= 3'b111;
      // memory_array[24047] <= 3'b111;
      // memory_array[24048] <= 3'b111;
      // memory_array[24049] <= 3'b101;
      // memory_array[24050] <= 3'b000;
      // memory_array[24051] <= 3'b000;
      // memory_array[24052] <= 3'b000;
      // memory_array[24053] <= 3'b000;
      // memory_array[24054] <= 3'b000;
      // memory_array[24055] <= 3'b000;
      // memory_array[24056] <= 3'b000;
      // memory_array[24057] <= 3'b000;
      // memory_array[24058] <= 3'b000;
      // memory_array[24059] <= 3'b000;
      // memory_array[24060] <= 3'b000;
      // memory_array[24061] <= 3'b000;
      // memory_array[24062] <= 3'b000;
      // memory_array[24063] <= 3'b000;
      // memory_array[24064] <= 3'b000;
      // memory_array[24065] <= 3'b000;
      // memory_array[24066] <= 3'b000;
      // memory_array[24067] <= 3'b000;
      // memory_array[24068] <= 3'b000;
      // memory_array[24069] <= 3'b000;
      // memory_array[24070] <= 3'b000;
      // memory_array[24071] <= 3'b000;
      // memory_array[24072] <= 3'b000;
      // memory_array[24073] <= 3'b101;
      // memory_array[24074] <= 3'b101;
      // memory_array[24075] <= 3'b000;
      // memory_array[24076] <= 3'b000;
      // memory_array[24077] <= 3'b000;
      // memory_array[24078] <= 3'b101;
      // memory_array[24079] <= 3'b000;
      // memory_array[24080] <= 3'b000;
      // memory_array[24081] <= 3'b000;
      // memory_array[24082] <= 3'b000;
      // memory_array[24083] <= 3'b000;
      // memory_array[24084] <= 3'b101;
      // memory_array[24085] <= 3'b000;
      // memory_array[24086] <= 3'b000;
      // memory_array[24087] <= 3'b000;
      // memory_array[24088] <= 3'b000;
      // memory_array[24089] <= 3'b000;
      // memory_array[24090] <= 3'b000;
      // memory_array[24091] <= 3'b000;
      // memory_array[24092] <= 3'b000;
      // memory_array[24093] <= 3'b000;
      // memory_array[24094] <= 3'b000;
      // memory_array[24095] <= 3'b000;
      // memory_array[24096] <= 3'b000;
      // memory_array[24097] <= 3'b000;
      // memory_array[24098] <= 3'b101;
      // memory_array[24099] <= 3'b101;
      // memory_array[24100] <= 3'b000;
      // memory_array[24101] <= 3'b000;
      // memory_array[24102] <= 3'b000;
      // memory_array[24103] <= 3'b000;
      // memory_array[24104] <= 3'b000;
      // memory_array[24105] <= 3'b000;
      // memory_array[24106] <= 3'b101;
      // memory_array[24107] <= 3'b000;
      // memory_array[24108] <= 3'b000;
      // memory_array[24109] <= 3'b101;
      // memory_array[24110] <= 3'b101;
      // memory_array[24111] <= 3'b101;
      // memory_array[24112] <= 3'b101;
      // memory_array[24113] <= 3'b101;
      // memory_array[24114] <= 3'b000;
      // memory_array[24115] <= 3'b000;
      // memory_array[24116] <= 3'b000;
      // memory_array[24117] <= 3'b000;
      // memory_array[24118] <= 3'b000;
      // memory_array[24119] <= 3'b000;
      // memory_array[24120] <= 3'b000;
      // memory_array[24121] <= 3'b000;
      // memory_array[24122] <= 3'b000;
      // memory_array[24123] <= 3'b000;
      // memory_array[24124] <= 3'b000;
      // memory_array[24125] <= 3'b000;
      // memory_array[24126] <= 3'b000;
      // memory_array[24127] <= 3'b000;
      // memory_array[24128] <= 3'b000;
      // memory_array[24129] <= 3'b000;
      // memory_array[24130] <= 3'b000;
      // memory_array[24131] <= 3'b000;
      // memory_array[24132] <= 3'b000;
      // memory_array[24133] <= 3'b000;
      // memory_array[24134] <= 3'b000;
      // memory_array[24135] <= 3'b000;
      // memory_array[24136] <= 3'b000;
      // memory_array[24137] <= 3'b000;
      // memory_array[24138] <= 3'b000;
      // memory_array[24139] <= 3'b000;
      // memory_array[24140] <= 3'b000;
      // memory_array[24141] <= 3'b000;
      // memory_array[24142] <= 3'b000;
      // memory_array[24143] <= 3'b101;
      // memory_array[24144] <= 3'b101;
      // memory_array[24145] <= 3'b000;
      // memory_array[24146] <= 3'b000;
      // memory_array[24147] <= 3'b000;
      // memory_array[24148] <= 3'b101;
      // memory_array[24149] <= 3'b000;
      // memory_array[24150] <= 3'b111;
      // memory_array[24151] <= 3'b111;
      // memory_array[24152] <= 3'b111;
      // memory_array[24153] <= 3'b111;
      // memory_array[24154] <= 3'b111;
      // memory_array[24155] <= 3'b101;
      // memory_array[24156] <= 3'b110;
      // memory_array[24157] <= 3'b000;
      // memory_array[24158] <= 3'b110;
      // memory_array[24159] <= 3'b110;
      // memory_array[24160] <= 3'b000;
      // memory_array[24161] <= 3'b000;
      // memory_array[24162] <= 3'b000;
      // memory_array[24163] <= 3'b000;
      // memory_array[24164] <= 3'b111;
      // memory_array[24165] <= 3'b111;
      // memory_array[24166] <= 3'b111;
      // memory_array[24167] <= 3'b000;
      // memory_array[24168] <= 3'b000;
      // memory_array[24169] <= 3'b111;
      // memory_array[24170] <= 3'b111;
      // memory_array[24171] <= 3'b111;
      // memory_array[24172] <= 3'b111;
      // memory_array[24173] <= 3'b111;
      // memory_array[24174] <= 3'b111;
      // memory_array[24175] <= 3'b111;
      // memory_array[24176] <= 3'b111;
      // memory_array[24177] <= 3'b111;
      // memory_array[24178] <= 3'b111;
      // memory_array[24179] <= 3'b110;
      // memory_array[24180] <= 3'b111;
      // memory_array[24181] <= 3'b111;
      // memory_array[24182] <= 3'b111;
      // memory_array[24183] <= 3'b110;
      // memory_array[24184] <= 3'b110;
      // memory_array[24185] <= 3'b111;
      // memory_array[24186] <= 3'b111;
      // memory_array[24187] <= 3'b111;
      // memory_array[24188] <= 3'b110;
      // memory_array[24189] <= 3'b000;
      // memory_array[24190] <= 3'b000;
      // memory_array[24191] <= 3'b101;
      // memory_array[24192] <= 3'b000;
      // memory_array[24193] <= 3'b110;
      // memory_array[24194] <= 3'b110;
      // memory_array[24195] <= 3'b000;
      // memory_array[24196] <= 3'b000;
      // memory_array[24197] <= 3'b000;
      // memory_array[24198] <= 3'b110;
      // memory_array[24199] <= 3'b110;
      // memory_array[24200] <= 3'b101;
      // memory_array[24201] <= 3'b110;
      // memory_array[24202] <= 3'b110;
      // memory_array[24203] <= 3'b000;
      // memory_array[24204] <= 3'b000;
      // memory_array[24205] <= 3'b110;
      // memory_array[24206] <= 3'b110;
      // memory_array[24207] <= 3'b101;
      // memory_array[24208] <= 3'b101;
      // memory_array[24209] <= 3'b000;
      // memory_array[24210] <= 3'b000;
      // memory_array[24211] <= 3'b110;
      // memory_array[24212] <= 3'b110;
      // memory_array[24213] <= 3'b110;
      // memory_array[24214] <= 3'b110;
      // memory_array[24215] <= 3'b110;
      // memory_array[24216] <= 3'b110;
      // memory_array[24217] <= 3'b110;
      // memory_array[24218] <= 3'b000;
      // memory_array[24219] <= 3'b000;
      // memory_array[24220] <= 3'b110;
      // memory_array[24221] <= 3'b000;
      // memory_array[24222] <= 3'b110;
      // memory_array[24223] <= 3'b000;
      // memory_array[24224] <= 3'b111;
      // memory_array[24225] <= 3'b111;
      // memory_array[24226] <= 3'b111;
      // memory_array[24227] <= 3'b000;
      // memory_array[24228] <= 3'b000;
      // memory_array[24229] <= 3'b000;
      // memory_array[24230] <= 3'b110;
      // memory_array[24231] <= 3'b110;
      // memory_array[24232] <= 3'b000;
      // memory_array[24233] <= 3'b111;
      // memory_array[24234] <= 3'b111;
      // memory_array[24235] <= 3'b111;
      // memory_array[24236] <= 3'b000;
      // memory_array[24237] <= 3'b110;
      // memory_array[24238] <= 3'b000;
      // memory_array[24239] <= 3'b000;
      // memory_array[24240] <= 3'b110;
      // memory_array[24241] <= 3'b110;
      // memory_array[24242] <= 3'b110;
      // memory_array[24243] <= 3'b000;
      // memory_array[24244] <= 3'b111;
      // memory_array[24245] <= 3'b111;
      // memory_array[24246] <= 3'b111;
      // memory_array[24247] <= 3'b111;
      // memory_array[24248] <= 3'b111;
      // memory_array[24249] <= 3'b101;
      // memory_array[24250] <= 3'b000;
      // memory_array[24251] <= 3'b000;
      // memory_array[24252] <= 3'b000;
      // memory_array[24253] <= 3'b000;
      // memory_array[24254] <= 3'b000;
      // memory_array[24255] <= 3'b000;
      // memory_array[24256] <= 3'b000;
      // memory_array[24257] <= 3'b000;
      // memory_array[24258] <= 3'b000;
      // memory_array[24259] <= 3'b000;
      // memory_array[24260] <= 3'b000;
      // memory_array[24261] <= 3'b000;
      // memory_array[24262] <= 3'b000;
      // memory_array[24263] <= 3'b000;
      // memory_array[24264] <= 3'b000;
      // memory_array[24265] <= 3'b101;
      // memory_array[24266] <= 3'b101;
      // memory_array[24267] <= 3'b000;
      // memory_array[24268] <= 3'b000;
      // memory_array[24269] <= 3'b000;
      // memory_array[24270] <= 3'b101;
      // memory_array[24271] <= 3'b101;
      // memory_array[24272] <= 3'b101;
      // memory_array[24273] <= 3'b000;
      // memory_array[24274] <= 3'b000;
      // memory_array[24275] <= 3'b101;
      // memory_array[24276] <= 3'b000;
      // memory_array[24277] <= 3'b000;
      // memory_array[24278] <= 3'b000;
      // memory_array[24279] <= 3'b000;
      // memory_array[24280] <= 3'b000;
      // memory_array[24281] <= 3'b101;
      // memory_array[24282] <= 3'b000;
      // memory_array[24283] <= 3'b000;
      // memory_array[24284] <= 3'b000;
      // memory_array[24285] <= 3'b000;
      // memory_array[24286] <= 3'b000;
      // memory_array[24287] <= 3'b000;
      // memory_array[24288] <= 3'b000;
      // memory_array[24289] <= 3'b000;
      // memory_array[24290] <= 3'b000;
      // memory_array[24291] <= 3'b000;
      // memory_array[24292] <= 3'b000;
      // memory_array[24293] <= 3'b000;
      // memory_array[24294] <= 3'b000;
      // memory_array[24295] <= 3'b101;
      // memory_array[24296] <= 3'b101;
      // memory_array[24297] <= 3'b101;
      // memory_array[24298] <= 3'b000;
      // memory_array[24299] <= 3'b000;
      // memory_array[24300] <= 3'b000;
      // memory_array[24301] <= 3'b101;
      // memory_array[24302] <= 3'b101;
      // memory_array[24303] <= 3'b000;
      // memory_array[24304] <= 3'b000;
      // memory_array[24305] <= 3'b000;
      // memory_array[24306] <= 3'b101;
      // memory_array[24307] <= 3'b101;
      // memory_array[24308] <= 3'b000;
      // memory_array[24309] <= 3'b101;
      // memory_array[24310] <= 3'b101;
      // memory_array[24311] <= 3'b101;
      // memory_array[24312] <= 3'b000;
      // memory_array[24313] <= 3'b000;
      // memory_array[24314] <= 3'b000;
      // memory_array[24315] <= 3'b000;
      // memory_array[24316] <= 3'b101;
      // memory_array[24317] <= 3'b000;
      // memory_array[24318] <= 3'b000;
      // memory_array[24319] <= 3'b000;
      // memory_array[24320] <= 3'b000;
      // memory_array[24321] <= 3'b101;
      // memory_array[24322] <= 3'b000;
      // memory_array[24323] <= 3'b000;
      // memory_array[24324] <= 3'b000;
      // memory_array[24325] <= 3'b000;
      // memory_array[24326] <= 3'b000;
      // memory_array[24327] <= 3'b000;
      // memory_array[24328] <= 3'b000;
      // memory_array[24329] <= 3'b000;
      // memory_array[24330] <= 3'b000;
      // memory_array[24331] <= 3'b000;
      // memory_array[24332] <= 3'b000;
      // memory_array[24333] <= 3'b000;
      // memory_array[24334] <= 3'b000;
      // memory_array[24335] <= 3'b000;
      // memory_array[24336] <= 3'b000;
      // memory_array[24337] <= 3'b000;
      // memory_array[24338] <= 3'b000;
      // memory_array[24339] <= 3'b000;
      // memory_array[24340] <= 3'b000;
      // memory_array[24341] <= 3'b000;
      // memory_array[24342] <= 3'b000;
      // memory_array[24343] <= 3'b000;
      // memory_array[24344] <= 3'b000;
      // memory_array[24345] <= 3'b101;
      // memory_array[24346] <= 3'b101;
      // memory_array[24347] <= 3'b000;
      // memory_array[24348] <= 3'b000;
      // memory_array[24349] <= 3'b000;
      // memory_array[24350] <= 3'b111;
      // memory_array[24351] <= 3'b111;
      // memory_array[24352] <= 3'b111;
      // memory_array[24353] <= 3'b111;
      // memory_array[24354] <= 3'b111;
      // memory_array[24355] <= 3'b101;
      // memory_array[24356] <= 3'b110;
      // memory_array[24357] <= 3'b110;
      // memory_array[24358] <= 3'b000;
      // memory_array[24359] <= 3'b000;
      // memory_array[24360] <= 3'b110;
      // memory_array[24361] <= 3'b000;
      // memory_array[24362] <= 3'b110;
      // memory_array[24363] <= 3'b000;
      // memory_array[24364] <= 3'b000;
      // memory_array[24365] <= 3'b000;
      // memory_array[24366] <= 3'b111;
      // memory_array[24367] <= 3'b111;
      // memory_array[24368] <= 3'b111;
      // memory_array[24369] <= 3'b000;
      // memory_array[24370] <= 3'b111;
      // memory_array[24371] <= 3'b111;
      // memory_array[24372] <= 3'b111;
      // memory_array[24373] <= 3'b111;
      // memory_array[24374] <= 3'b000;
      // memory_array[24375] <= 3'b111;
      // memory_array[24376] <= 3'b111;
      // memory_array[24377] <= 3'b111;
      // memory_array[24378] <= 3'b111;
      // memory_array[24379] <= 3'b111;
      // memory_array[24380] <= 3'b110;
      // memory_array[24381] <= 3'b110;
      // memory_array[24382] <= 3'b110;
      // memory_array[24383] <= 3'b000;
      // memory_array[24384] <= 3'b111;
      // memory_array[24385] <= 3'b110;
      // memory_array[24386] <= 3'b110;
      // memory_array[24387] <= 3'b110;
      // memory_array[24388] <= 3'b000;
      // memory_array[24389] <= 3'b000;
      // memory_array[24390] <= 3'b000;
      // memory_array[24391] <= 3'b101;
      // memory_array[24392] <= 3'b110;
      // memory_array[24393] <= 3'b000;
      // memory_array[24394] <= 3'b000;
      // memory_array[24395] <= 3'b110;
      // memory_array[24396] <= 3'b110;
      // memory_array[24397] <= 3'b110;
      // memory_array[24398] <= 3'b000;
      // memory_array[24399] <= 3'b101;
      // memory_array[24400] <= 3'b101;
      // memory_array[24401] <= 3'b101;
      // memory_array[24402] <= 3'b110;
      // memory_array[24403] <= 3'b101;
      // memory_array[24404] <= 3'b101;
      // memory_array[24405] <= 3'b110;
      // memory_array[24406] <= 3'b101;
      // memory_array[24407] <= 3'b101;
      // memory_array[24408] <= 3'b101;
      // memory_array[24409] <= 3'b000;
      // memory_array[24410] <= 3'b000;
      // memory_array[24411] <= 3'b110;
      // memory_array[24412] <= 3'b110;
      // memory_array[24413] <= 3'b110;
      // memory_array[24414] <= 3'b110;
      // memory_array[24415] <= 3'b110;
      // memory_array[24416] <= 3'b110;
      // memory_array[24417] <= 3'b110;
      // memory_array[24418] <= 3'b110;
      // memory_array[24419] <= 3'b110;
      // memory_array[24420] <= 3'b110;
      // memory_array[24421] <= 3'b000;
      // memory_array[24422] <= 3'b110;
      // memory_array[24423] <= 3'b000;
      // memory_array[24424] <= 3'b111;
      // memory_array[24425] <= 3'b111;
      // memory_array[24426] <= 3'b111;
      // memory_array[24427] <= 3'b111;
      // memory_array[24428] <= 3'b111;
      // memory_array[24429] <= 3'b111;
      // memory_array[24430] <= 3'b111;
      // memory_array[24431] <= 3'b111;
      // memory_array[24432] <= 3'b000;
      // memory_array[24433] <= 3'b110;
      // memory_array[24434] <= 3'b111;
      // memory_array[24435] <= 3'b110;
      // memory_array[24436] <= 3'b110;
      // memory_array[24437] <= 3'b110;
      // memory_array[24438] <= 3'b000;
      // memory_array[24439] <= 3'b111;
      // memory_array[24440] <= 3'b111;
      // memory_array[24441] <= 3'b111;
      // memory_array[24442] <= 3'b111;
      // memory_array[24443] <= 3'b111;
      // memory_array[24444] <= 3'b111;
      // memory_array[24445] <= 3'b111;
      // memory_array[24446] <= 3'b111;
      // memory_array[24447] <= 3'b111;
      // memory_array[24448] <= 3'b111;
      // memory_array[24449] <= 3'b111;
      // memory_array[24450] <= 3'b111;
      // memory_array[24451] <= 3'b111;
      // memory_array[24452] <= 3'b111;
      // memory_array[24453] <= 3'b111;
      // memory_array[24454] <= 3'b101;
      // memory_array[24455] <= 3'b000;
      // memory_array[24456] <= 3'b000;
      // memory_array[24457] <= 3'b000;
      // memory_array[24458] <= 3'b000;
      // memory_array[24459] <= 3'b000;
      // memory_array[24460] <= 3'b000;
      // memory_array[24461] <= 3'b000;
      // memory_array[24462] <= 3'b000;
      // memory_array[24463] <= 3'b000;
      // memory_array[24464] <= 3'b000;
      // memory_array[24465] <= 3'b101;
      // memory_array[24466] <= 3'b101;
      // memory_array[24467] <= 3'b101;
      // memory_array[24468] <= 3'b000;
      // memory_array[24469] <= 3'b000;
      // memory_array[24470] <= 3'b000;
      // memory_array[24471] <= 3'b000;
      // memory_array[24472] <= 3'b000;
      // memory_array[24473] <= 3'b000;
      // memory_array[24474] <= 3'b000;
      // memory_array[24475] <= 3'b101;
      // memory_array[24476] <= 3'b101;
      // memory_array[24477] <= 3'b101;
      // memory_array[24478] <= 3'b101;
      // memory_array[24479] <= 3'b000;
      // memory_array[24480] <= 3'b101;
      // memory_array[24481] <= 3'b000;
      // memory_array[24482] <= 3'b101;
      // memory_array[24483] <= 3'b000;
      // memory_array[24484] <= 3'b000;
      // memory_array[24485] <= 3'b000;
      // memory_array[24486] <= 3'b000;
      // memory_array[24487] <= 3'b110;
      // memory_array[24488] <= 3'b000;
      // memory_array[24489] <= 3'b000;
      // memory_array[24490] <= 3'b000;
      // memory_array[24491] <= 3'b000;
      // memory_array[24492] <= 3'b110;
      // memory_array[24493] <= 3'b000;
      // memory_array[24494] <= 3'b000;
      // memory_array[24495] <= 3'b101;
      // memory_array[24496] <= 3'b101;
      // memory_array[24497] <= 3'b101;
      // memory_array[24498] <= 3'b000;
      // memory_array[24499] <= 3'b000;
      // memory_array[24500] <= 3'b101;
      // memory_array[24501] <= 3'b101;
      // memory_array[24502] <= 3'b101;
      // memory_array[24503] <= 3'b000;
      // memory_array[24504] <= 3'b000;
      // memory_array[24505] <= 3'b000;
      // memory_array[24506] <= 3'b000;
      // memory_array[24507] <= 3'b000;
      // memory_array[24508] <= 3'b101;
      // memory_array[24509] <= 3'b000;
      // memory_array[24510] <= 3'b101;
      // memory_array[24511] <= 3'b101;
      // memory_array[24512] <= 3'b000;
      // memory_array[24513] <= 3'b000;
      // memory_array[24514] <= 3'b000;
      // memory_array[24515] <= 3'b000;
      // memory_array[24516] <= 3'b101;
      // memory_array[24517] <= 3'b000;
      // memory_array[24518] <= 3'b000;
      // memory_array[24519] <= 3'b101;
      // memory_array[24520] <= 3'b000;
      // memory_array[24521] <= 3'b000;
      // memory_array[24522] <= 3'b101;
      // memory_array[24523] <= 3'b000;
      // memory_array[24524] <= 3'b000;
      // memory_array[24525] <= 3'b000;
      // memory_array[24526] <= 3'b000;
      // memory_array[24527] <= 3'b101;
      // memory_array[24528] <= 3'b000;
      // memory_array[24529] <= 3'b000;
      // memory_array[24530] <= 3'b000;
      // memory_array[24531] <= 3'b000;
      // memory_array[24532] <= 3'b000;
      // memory_array[24533] <= 3'b000;
      // memory_array[24534] <= 3'b000;
      // memory_array[24535] <= 3'b101;
      // memory_array[24536] <= 3'b101;
      // memory_array[24537] <= 3'b101;
      // memory_array[24538] <= 3'b000;
      // memory_array[24539] <= 3'b000;
      // memory_array[24540] <= 3'b101;
      // memory_array[24541] <= 3'b101;
      // memory_array[24542] <= 3'b000;
      // memory_array[24543] <= 3'b000;
      // memory_array[24544] <= 3'b000;
      // memory_array[24545] <= 3'b111;
      // memory_array[24546] <= 3'b111;
      // memory_array[24547] <= 3'b111;
      // memory_array[24548] <= 3'b111;
      // memory_array[24549] <= 3'b111;
      // memory_array[24550] <= 3'b111;
      // memory_array[24551] <= 3'b111;
      // memory_array[24552] <= 3'b111;
      // memory_array[24553] <= 3'b111;
      // memory_array[24554] <= 3'b111;
      // memory_array[24555] <= 3'b111;
      // memory_array[24556] <= 3'b111;
      // memory_array[24557] <= 3'b111;
      // memory_array[24558] <= 3'b111;
      // memory_array[24559] <= 3'b111;
      // memory_array[24560] <= 3'b111;
      // memory_array[24561] <= 3'b000;
      // memory_array[24562] <= 3'b110;
      // memory_array[24563] <= 3'b110;
      // memory_array[24564] <= 3'b110;
      // memory_array[24565] <= 3'b110;
      // memory_array[24566] <= 3'b110;
      // memory_array[24567] <= 3'b110;
      // memory_array[24568] <= 3'b111;
      // memory_array[24569] <= 3'b111;
      // memory_array[24570] <= 3'b000;
      // memory_array[24571] <= 3'b000;
      // memory_array[24572] <= 3'b000;
      // memory_array[24573] <= 3'b000;
      // memory_array[24574] <= 3'b111;
      // memory_array[24575] <= 3'b111;
      // memory_array[24576] <= 3'b111;
      // memory_array[24577] <= 3'b111;
      // memory_array[24578] <= 3'b111;
      // memory_array[24579] <= 3'b111;
      // memory_array[24580] <= 3'b110;
      // memory_array[24581] <= 3'b110;
      // memory_array[24582] <= 3'b110;
      // memory_array[24583] <= 3'b110;
      // memory_array[24584] <= 3'b000;
      // memory_array[24585] <= 3'b110;
      // memory_array[24586] <= 3'b110;
      // memory_array[24587] <= 3'b110;
      // memory_array[24588] <= 3'b000;
      // memory_array[24589] <= 3'b000;
      // memory_array[24590] <= 3'b000;
      // memory_array[24591] <= 3'b101;
      // memory_array[24592] <= 3'b101;
      // memory_array[24593] <= 3'b101;
      // memory_array[24594] <= 3'b000;
      // memory_array[24595] <= 3'b101;
      // memory_array[24596] <= 3'b101;
      // memory_array[24597] <= 3'b110;
      // memory_array[24598] <= 3'b101;
      // memory_array[24599] <= 3'b101;
      // memory_array[24600] <= 3'b101;
      // memory_array[24601] <= 3'b101;
      // memory_array[24602] <= 3'b101;
      // memory_array[24603] <= 3'b111;
      // memory_array[24604] <= 3'b111;
      // memory_array[24605] <= 3'b101;
      // memory_array[24606] <= 3'b101;
      // memory_array[24607] <= 3'b101;
      // memory_array[24608] <= 3'b101;
      // memory_array[24609] <= 3'b000;
      // memory_array[24610] <= 3'b000;
      // memory_array[24611] <= 3'b110;
      // memory_array[24612] <= 3'b000;
      // memory_array[24613] <= 3'b110;
      // memory_array[24614] <= 3'b110;
      // memory_array[24615] <= 3'b000;
      // memory_array[24616] <= 3'b110;
      // memory_array[24617] <= 3'b111;
      // memory_array[24618] <= 3'b110;
      // memory_array[24619] <= 3'b110;
      // memory_array[24620] <= 3'b111;
      // memory_array[24621] <= 3'b000;
      // memory_array[24622] <= 3'b110;
      // memory_array[24623] <= 3'b000;
      // memory_array[24624] <= 3'b111;
      // memory_array[24625] <= 3'b111;
      // memory_array[24626] <= 3'b111;
      // memory_array[24627] <= 3'b111;
      // memory_array[24628] <= 3'b111;
      // memory_array[24629] <= 3'b111;
      // memory_array[24630] <= 3'b000;
      // memory_array[24631] <= 3'b000;
      // memory_array[24632] <= 3'b000;
      // memory_array[24633] <= 3'b110;
      // memory_array[24634] <= 3'b110;
      // memory_array[24635] <= 3'b110;
      // memory_array[24636] <= 3'b110;
      // memory_array[24637] <= 3'b110;
      // memory_array[24638] <= 3'b000;
      // memory_array[24639] <= 3'b111;
      // memory_array[24640] <= 3'b111;
      // memory_array[24641] <= 3'b111;
      // memory_array[24642] <= 3'b111;
      // memory_array[24643] <= 3'b111;
      // memory_array[24644] <= 3'b111;
      // memory_array[24645] <= 3'b111;
      // memory_array[24646] <= 3'b111;
      // memory_array[24647] <= 3'b111;
      // memory_array[24648] <= 3'b111;
      // memory_array[24649] <= 3'b111;
      // memory_array[24650] <= 3'b111;
      // memory_array[24651] <= 3'b111;
      // memory_array[24652] <= 3'b111;
      // memory_array[24653] <= 3'b111;
      // memory_array[24654] <= 3'b101;
      // memory_array[24655] <= 3'b000;
      // memory_array[24656] <= 3'b000;
      // memory_array[24657] <= 3'b000;
      // memory_array[24658] <= 3'b000;
      // memory_array[24659] <= 3'b000;
      // memory_array[24660] <= 3'b000;
      // memory_array[24661] <= 3'b000;
      // memory_array[24662] <= 3'b000;
      // memory_array[24663] <= 3'b101;
      // memory_array[24664] <= 3'b101;
      // memory_array[24665] <= 3'b000;
      // memory_array[24666] <= 3'b000;
      // memory_array[24667] <= 3'b000;
      // memory_array[24668] <= 3'b000;
      // memory_array[24669] <= 3'b000;
      // memory_array[24670] <= 3'b000;
      // memory_array[24671] <= 3'b000;
      // memory_array[24672] <= 3'b000;
      // memory_array[24673] <= 3'b101;
      // memory_array[24674] <= 3'b101;
      // memory_array[24675] <= 3'b000;
      // memory_array[24676] <= 3'b000;
      // memory_array[24677] <= 3'b000;
      // memory_array[24678] <= 3'b101;
      // memory_array[24679] <= 3'b000;
      // memory_array[24680] <= 3'b000;
      // memory_array[24681] <= 3'b000;
      // memory_array[24682] <= 3'b101;
      // memory_array[24683] <= 3'b101;
      // memory_array[24684] <= 3'b000;
      // memory_array[24685] <= 3'b000;
      // memory_array[24686] <= 3'b000;
      // memory_array[24687] <= 3'b000;
      // memory_array[24688] <= 3'b000;
      // memory_array[24689] <= 3'b000;
      // memory_array[24690] <= 3'b000;
      // memory_array[24691] <= 3'b000;
      // memory_array[24692] <= 3'b000;
      // memory_array[24693] <= 3'b110;
      // memory_array[24694] <= 3'b101;
      // memory_array[24695] <= 3'b000;
      // memory_array[24696] <= 3'b000;
      // memory_array[24697] <= 3'b000;
      // memory_array[24698] <= 3'b101;
      // memory_array[24699] <= 3'b101;
      // memory_array[24700] <= 3'b000;
      // memory_array[24701] <= 3'b000;
      // memory_array[24702] <= 3'b000;
      // memory_array[24703] <= 3'b101;
      // memory_array[24704] <= 3'b101;
      // memory_array[24705] <= 3'b000;
      // memory_array[24706] <= 3'b000;
      // memory_array[24707] <= 3'b000;
      // memory_array[24708] <= 3'b000;
      // memory_array[24709] <= 3'b000;
      // memory_array[24710] <= 3'b000;
      // memory_array[24711] <= 3'b101;
      // memory_array[24712] <= 3'b101;
      // memory_array[24713] <= 3'b000;
      // memory_array[24714] <= 3'b101;
      // memory_array[24715] <= 3'b101;
      // memory_array[24716] <= 3'b000;
      // memory_array[24717] <= 3'b000;
      // memory_array[24718] <= 3'b000;
      // memory_array[24719] <= 3'b000;
      // memory_array[24720] <= 3'b000;
      // memory_array[24721] <= 3'b101;
      // memory_array[24722] <= 3'b000;
      // memory_array[24723] <= 3'b000;
      // memory_array[24724] <= 3'b101;
      // memory_array[24725] <= 3'b000;
      // memory_array[24726] <= 3'b000;
      // memory_array[24727] <= 3'b000;
      // memory_array[24728] <= 3'b000;
      // memory_array[24729] <= 3'b101;
      // memory_array[24730] <= 3'b000;
      // memory_array[24731] <= 3'b000;
      // memory_array[24732] <= 3'b000;
      // memory_array[24733] <= 3'b000;
      // memory_array[24734] <= 3'b101;
      // memory_array[24735] <= 3'b000;
      // memory_array[24736] <= 3'b000;
      // memory_array[24737] <= 3'b000;
      // memory_array[24738] <= 3'b000;
      // memory_array[24739] <= 3'b000;
      // memory_array[24740] <= 3'b000;
      // memory_array[24741] <= 3'b000;
      // memory_array[24742] <= 3'b000;
      // memory_array[24743] <= 3'b000;
      // memory_array[24744] <= 3'b000;
      // memory_array[24745] <= 3'b111;
      // memory_array[24746] <= 3'b111;
      // memory_array[24747] <= 3'b111;
      // memory_array[24748] <= 3'b111;
      // memory_array[24749] <= 3'b111;
      // memory_array[24750] <= 3'b111;
      // memory_array[24751] <= 3'b111;
      // memory_array[24752] <= 3'b111;
      // memory_array[24753] <= 3'b111;
      // memory_array[24754] <= 3'b111;
      // memory_array[24755] <= 3'b111;
      // memory_array[24756] <= 3'b111;
      // memory_array[24757] <= 3'b111;
      // memory_array[24758] <= 3'b111;
      // memory_array[24759] <= 3'b111;
      // memory_array[24760] <= 3'b111;
      // memory_array[24761] <= 3'b000;
      // memory_array[24762] <= 3'b111;
      // memory_array[24763] <= 3'b110;
      // memory_array[24764] <= 3'b110;
      // memory_array[24765] <= 3'b111;
      // memory_array[24766] <= 3'b110;
      // memory_array[24767] <= 3'b111;
      // memory_array[24768] <= 3'b110;
      // memory_array[24769] <= 3'b110;
      // memory_array[24770] <= 3'b110;
      // memory_array[24771] <= 3'b110;
      // memory_array[24772] <= 3'b000;
      // memory_array[24773] <= 3'b111;
      // memory_array[24774] <= 3'b111;
      // memory_array[24775] <= 3'b111;
      // memory_array[24776] <= 3'b111;
      // memory_array[24777] <= 3'b111;
      // memory_array[24778] <= 3'b111;
      // memory_array[24779] <= 3'b110;
      // memory_array[24780] <= 3'b110;
      // memory_array[24781] <= 3'b110;
      // memory_array[24782] <= 3'b110;
      // memory_array[24783] <= 3'b110;
      // memory_array[24784] <= 3'b110;
      // memory_array[24785] <= 3'b000;
      // memory_array[24786] <= 3'b000;
      // memory_array[24787] <= 3'b000;
      // memory_array[24788] <= 3'b110;
      // memory_array[24789] <= 3'b000;
      // memory_array[24790] <= 3'b000;
      // memory_array[24791] <= 3'b101;
      // memory_array[24792] <= 3'b101;
      // memory_array[24793] <= 3'b101;
      // memory_array[24794] <= 3'b101;
      // memory_array[24795] <= 3'b111;
      // memory_array[24796] <= 3'b111;
      // memory_array[24797] <= 3'b101;
      // memory_array[24798] <= 3'b101;
      // memory_array[24799] <= 3'b101;
      // memory_array[24800] <= 3'b101;
      // memory_array[24801] <= 3'b101;
      // memory_array[24802] <= 3'b101;
      // memory_array[24803] <= 3'b101;
      // memory_array[24804] <= 3'b101;
      // memory_array[24805] <= 3'b101;
      // memory_array[24806] <= 3'b101;
      // memory_array[24807] <= 3'b101;
      // memory_array[24808] <= 3'b101;
      // memory_array[24809] <= 3'b000;
      // memory_array[24810] <= 3'b000;
      // memory_array[24811] <= 3'b110;
      // memory_array[24812] <= 3'b000;
      // memory_array[24813] <= 3'b110;
      // memory_array[24814] <= 3'b110;
      // memory_array[24815] <= 3'b000;
      // memory_array[24816] <= 3'b110;
      // memory_array[24817] <= 3'b111;
      // memory_array[24818] <= 3'b110;
      // memory_array[24819] <= 3'b110;
      // memory_array[24820] <= 3'b111;
      // memory_array[24821] <= 3'b000;
      // memory_array[24822] <= 3'b000;
      // memory_array[24823] <= 3'b111;
      // memory_array[24824] <= 3'b111;
      // memory_array[24825] <= 3'b111;
      // memory_array[24826] <= 3'b111;
      // memory_array[24827] <= 3'b000;
      // memory_array[24828] <= 3'b000;
      // memory_array[24829] <= 3'b110;
      // memory_array[24830] <= 3'b111;
      // memory_array[24831] <= 3'b111;
      // memory_array[24832] <= 3'b000;
      // memory_array[24833] <= 3'b110;
      // memory_array[24834] <= 3'b110;
      // memory_array[24835] <= 3'b110;
      // memory_array[24836] <= 3'b110;
      // memory_array[24837] <= 3'b000;
      // memory_array[24838] <= 3'b000;
      // memory_array[24839] <= 3'b111;
      // memory_array[24840] <= 3'b111;
      // memory_array[24841] <= 3'b111;
      // memory_array[24842] <= 3'b111;
      // memory_array[24843] <= 3'b111;
      // memory_array[24844] <= 3'b111;
      // memory_array[24845] <= 3'b111;
      // memory_array[24846] <= 3'b111;
      // memory_array[24847] <= 3'b111;
      // memory_array[24848] <= 3'b111;
      // memory_array[24849] <= 3'b111;
      // memory_array[24850] <= 3'b111;
      // memory_array[24851] <= 3'b111;
      // memory_array[24852] <= 3'b111;
      // memory_array[24853] <= 3'b111;
      // memory_array[24854] <= 3'b101;
      // memory_array[24855] <= 3'b000;
      // memory_array[24856] <= 3'b000;
      // memory_array[24857] <= 3'b000;
      // memory_array[24858] <= 3'b000;
      // memory_array[24859] <= 3'b000;
      // memory_array[24860] <= 3'b000;
      // memory_array[24861] <= 3'b000;
      // memory_array[24862] <= 3'b000;
      // memory_array[24863] <= 3'b000;
      // memory_array[24864] <= 3'b000;
      // memory_array[24865] <= 3'b000;
      // memory_array[24866] <= 3'b000;
      // memory_array[24867] <= 3'b000;
      // memory_array[24868] <= 3'b000;
      // memory_array[24869] <= 3'b000;
      // memory_array[24870] <= 3'b000;
      // memory_array[24871] <= 3'b101;
      // memory_array[24872] <= 3'b000;
      // memory_array[24873] <= 3'b101;
      // memory_array[24874] <= 3'b000;
      // memory_array[24875] <= 3'b101;
      // memory_array[24876] <= 3'b000;
      // memory_array[24877] <= 3'b000;
      // memory_array[24878] <= 3'b000;
      // memory_array[24879] <= 3'b000;
      // memory_array[24880] <= 3'b000;
      // memory_array[24881] <= 3'b000;
      // memory_array[24882] <= 3'b000;
      // memory_array[24883] <= 3'b101;
      // memory_array[24884] <= 3'b000;
      // memory_array[24885] <= 3'b000;
      // memory_array[24886] <= 3'b000;
      // memory_array[24887] <= 3'b000;
      // memory_array[24888] <= 3'b110;
      // memory_array[24889] <= 3'b000;
      // memory_array[24890] <= 3'b000;
      // memory_array[24891] <= 3'b000;
      // memory_array[24892] <= 3'b000;
      // memory_array[24893] <= 3'b110;
      // memory_array[24894] <= 3'b101;
      // memory_array[24895] <= 3'b000;
      // memory_array[24896] <= 3'b000;
      // memory_array[24897] <= 3'b000;
      // memory_array[24898] <= 3'b101;
      // memory_array[24899] <= 3'b101;
      // memory_array[24900] <= 3'b000;
      // memory_array[24901] <= 3'b000;
      // memory_array[24902] <= 3'b000;
      // memory_array[24903] <= 3'b101;
      // memory_array[24904] <= 3'b101;
      // memory_array[24905] <= 3'b000;
      // memory_array[24906] <= 3'b000;
      // memory_array[24907] <= 3'b000;
      // memory_array[24908] <= 3'b000;
      // memory_array[24909] <= 3'b101;
      // memory_array[24910] <= 3'b101;
      // memory_array[24911] <= 3'b101;
      // memory_array[24912] <= 3'b000;
      // memory_array[24913] <= 3'b101;
      // memory_array[24914] <= 3'b000;
      // memory_array[24915] <= 3'b000;
      // memory_array[24916] <= 3'b000;
      // memory_array[24917] <= 3'b000;
      // memory_array[24918] <= 3'b000;
      // memory_array[24919] <= 3'b000;
      // memory_array[24920] <= 3'b000;
      // memory_array[24921] <= 3'b000;
      // memory_array[24922] <= 3'b000;
      // memory_array[24923] <= 3'b101;
      // memory_array[24924] <= 3'b000;
      // memory_array[24925] <= 3'b000;
      // memory_array[24926] <= 3'b000;
      // memory_array[24927] <= 3'b000;
      // memory_array[24928] <= 3'b000;
      // memory_array[24929] <= 3'b000;
      // memory_array[24930] <= 3'b000;
      // memory_array[24931] <= 3'b000;
      // memory_array[24932] <= 3'b000;
      // memory_array[24933] <= 3'b101;
      // memory_array[24934] <= 3'b101;
      // memory_array[24935] <= 3'b000;
      // memory_array[24936] <= 3'b000;
      // memory_array[24937] <= 3'b000;
      // memory_array[24938] <= 3'b101;
      // memory_array[24939] <= 3'b000;
      // memory_array[24940] <= 3'b000;
      // memory_array[24941] <= 3'b000;
      // memory_array[24942] <= 3'b000;
      // memory_array[24943] <= 3'b000;
      // memory_array[24944] <= 3'b000;
      // memory_array[24945] <= 3'b111;
      // memory_array[24946] <= 3'b111;
      // memory_array[24947] <= 3'b111;
      // memory_array[24948] <= 3'b111;
      // memory_array[24949] <= 3'b111;
      // memory_array[24950] <= 3'b111;
      // memory_array[24951] <= 3'b111;
      // memory_array[24952] <= 3'b111;
      // memory_array[24953] <= 3'b111;
      // memory_array[24954] <= 3'b111;
      // memory_array[24955] <= 3'b111;
      // memory_array[24956] <= 3'b111;
      // memory_array[24957] <= 3'b111;
      // memory_array[24958] <= 3'b111;
      // memory_array[24959] <= 3'b111;
      // memory_array[24960] <= 3'b111;
      // memory_array[24961] <= 3'b000;
      // memory_array[24962] <= 3'b111;
      // memory_array[24963] <= 3'b110;
      // memory_array[24964] <= 3'b110;
      // memory_array[24965] <= 3'b111;
      // memory_array[24966] <= 3'b110;
      // memory_array[24967] <= 3'b111;
      // memory_array[24968] <= 3'b110;
      // memory_array[24969] <= 3'b110;
      // memory_array[24970] <= 3'b110;
      // memory_array[24971] <= 3'b110;
      // memory_array[24972] <= 3'b000;
      // memory_array[24973] <= 3'b110;
      // memory_array[24974] <= 3'b000;
      // memory_array[24975] <= 3'b000;
      // memory_array[24976] <= 3'b111;
      // memory_array[24977] <= 3'b111;
      // memory_array[24978] <= 3'b111;
      // memory_array[24979] <= 3'b000;
      // memory_array[24980] <= 3'b110;
      // memory_array[24981] <= 3'b110;
      // memory_array[24982] <= 3'b110;
      // memory_array[24983] <= 3'b110;
      // memory_array[24984] <= 3'b110;
      // memory_array[24985] <= 3'b000;
      // memory_array[24986] <= 3'b000;
      // memory_array[24987] <= 3'b000;
      // memory_array[24988] <= 3'b110;
      // memory_array[24989] <= 3'b000;
      // memory_array[24990] <= 3'b000;
      // memory_array[24991] <= 3'b101;
      // memory_array[24992] <= 3'b111;
      // memory_array[24993] <= 3'b101;
      // memory_array[24994] <= 3'b101;
      // memory_array[24995] <= 3'b101;
      // memory_array[24996] <= 3'b101;
      // memory_array[24997] <= 3'b101;
      // memory_array[24998] <= 3'b101;
      // memory_array[24999] <= 3'b101;
      // memory_array[25000] <= 3'b101;
      // memory_array[25001] <= 3'b101;
      // memory_array[25002] <= 3'b101;
      // memory_array[25003] <= 3'b101;
      // memory_array[25004] <= 3'b101;
      // memory_array[25005] <= 3'b101;
      // memory_array[25006] <= 3'b101;
      // memory_array[25007] <= 3'b101;
      // memory_array[25008] <= 3'b101;
      // memory_array[25009] <= 3'b000;
      // memory_array[25010] <= 3'b000;
      // memory_array[25011] <= 3'b110;
      // memory_array[25012] <= 3'b000;
      // memory_array[25013] <= 3'b110;
      // memory_array[25014] <= 3'b110;
      // memory_array[25015] <= 3'b000;
      // memory_array[25016] <= 3'b110;
      // memory_array[25017] <= 3'b111;
      // memory_array[25018] <= 3'b110;
      // memory_array[25019] <= 3'b110;
      // memory_array[25020] <= 3'b111;
      // memory_array[25021] <= 3'b000;
      // memory_array[25022] <= 3'b000;
      // memory_array[25023] <= 3'b111;
      // memory_array[25024] <= 3'b111;
      // memory_array[25025] <= 3'b111;
      // memory_array[25026] <= 3'b111;
      // memory_array[25027] <= 3'b000;
      // memory_array[25028] <= 3'b000;
      // memory_array[25029] <= 3'b110;
      // memory_array[25030] <= 3'b111;
      // memory_array[25031] <= 3'b111;
      // memory_array[25032] <= 3'b000;
      // memory_array[25033] <= 3'b110;
      // memory_array[25034] <= 3'b110;
      // memory_array[25035] <= 3'b110;
      // memory_array[25036] <= 3'b110;
      // memory_array[25037] <= 3'b000;
      // memory_array[25038] <= 3'b000;
      // memory_array[25039] <= 3'b111;
      // memory_array[25040] <= 3'b111;
      // memory_array[25041] <= 3'b111;
      // memory_array[25042] <= 3'b111;
      // memory_array[25043] <= 3'b111;
      // memory_array[25044] <= 3'b111;
      // memory_array[25045] <= 3'b111;
      // memory_array[25046] <= 3'b111;
      // memory_array[25047] <= 3'b111;
      // memory_array[25048] <= 3'b111;
      // memory_array[25049] <= 3'b111;
      // memory_array[25050] <= 3'b111;
      // memory_array[25051] <= 3'b111;
      // memory_array[25052] <= 3'b111;
      // memory_array[25053] <= 3'b111;
      // memory_array[25054] <= 3'b101;
      // memory_array[25055] <= 3'b000;
      // memory_array[25056] <= 3'b000;
      // memory_array[25057] <= 3'b000;
      // memory_array[25058] <= 3'b000;
      // memory_array[25059] <= 3'b000;
      // memory_array[25060] <= 3'b000;
      // memory_array[25061] <= 3'b000;
      // memory_array[25062] <= 3'b000;
      // memory_array[25063] <= 3'b000;
      // memory_array[25064] <= 3'b000;
      // memory_array[25065] <= 3'b000;
      // memory_array[25066] <= 3'b000;
      // memory_array[25067] <= 3'b000;
      // memory_array[25068] <= 3'b000;
      // memory_array[25069] <= 3'b000;
      // memory_array[25070] <= 3'b000;
      // memory_array[25071] <= 3'b101;
      // memory_array[25072] <= 3'b000;
      // memory_array[25073] <= 3'b101;
      // memory_array[25074] <= 3'b000;
      // memory_array[25075] <= 3'b101;
      // memory_array[25076] <= 3'b000;
      // memory_array[25077] <= 3'b000;
      // memory_array[25078] <= 3'b000;
      // memory_array[25079] <= 3'b000;
      // memory_array[25080] <= 3'b000;
      // memory_array[25081] <= 3'b000;
      // memory_array[25082] <= 3'b000;
      // memory_array[25083] <= 3'b101;
      // memory_array[25084] <= 3'b000;
      // memory_array[25085] <= 3'b000;
      // memory_array[25086] <= 3'b000;
      // memory_array[25087] <= 3'b000;
      // memory_array[25088] <= 3'b110;
      // memory_array[25089] <= 3'b000;
      // memory_array[25090] <= 3'b000;
      // memory_array[25091] <= 3'b000;
      // memory_array[25092] <= 3'b000;
      // memory_array[25093] <= 3'b110;
      // memory_array[25094] <= 3'b101;
      // memory_array[25095] <= 3'b000;
      // memory_array[25096] <= 3'b000;
      // memory_array[25097] <= 3'b000;
      // memory_array[25098] <= 3'b101;
      // memory_array[25099] <= 3'b101;
      // memory_array[25100] <= 3'b000;
      // memory_array[25101] <= 3'b000;
      // memory_array[25102] <= 3'b000;
      // memory_array[25103] <= 3'b101;
      // memory_array[25104] <= 3'b101;
      // memory_array[25105] <= 3'b000;
      // memory_array[25106] <= 3'b000;
      // memory_array[25107] <= 3'b000;
      // memory_array[25108] <= 3'b000;
      // memory_array[25109] <= 3'b101;
      // memory_array[25110] <= 3'b101;
      // memory_array[25111] <= 3'b101;
      // memory_array[25112] <= 3'b000;
      // memory_array[25113] <= 3'b101;
      // memory_array[25114] <= 3'b000;
      // memory_array[25115] <= 3'b000;
      // memory_array[25116] <= 3'b000;
      // memory_array[25117] <= 3'b000;
      // memory_array[25118] <= 3'b000;
      // memory_array[25119] <= 3'b000;
      // memory_array[25120] <= 3'b000;
      // memory_array[25121] <= 3'b000;
      // memory_array[25122] <= 3'b000;
      // memory_array[25123] <= 3'b101;
      // memory_array[25124] <= 3'b000;
      // memory_array[25125] <= 3'b000;
      // memory_array[25126] <= 3'b000;
      // memory_array[25127] <= 3'b000;
      // memory_array[25128] <= 3'b000;
      // memory_array[25129] <= 3'b000;
      // memory_array[25130] <= 3'b000;
      // memory_array[25131] <= 3'b000;
      // memory_array[25132] <= 3'b000;
      // memory_array[25133] <= 3'b101;
      // memory_array[25134] <= 3'b101;
      // memory_array[25135] <= 3'b000;
      // memory_array[25136] <= 3'b000;
      // memory_array[25137] <= 3'b000;
      // memory_array[25138] <= 3'b101;
      // memory_array[25139] <= 3'b000;
      // memory_array[25140] <= 3'b000;
      // memory_array[25141] <= 3'b000;
      // memory_array[25142] <= 3'b000;
      // memory_array[25143] <= 3'b000;
      // memory_array[25144] <= 3'b000;
      // memory_array[25145] <= 3'b111;
      // memory_array[25146] <= 3'b111;
      // memory_array[25147] <= 3'b111;
      // memory_array[25148] <= 3'b111;
      // memory_array[25149] <= 3'b111;
      // memory_array[25150] <= 3'b111;
      // memory_array[25151] <= 3'b111;
      // memory_array[25152] <= 3'b111;
      // memory_array[25153] <= 3'b111;
      // memory_array[25154] <= 3'b111;
      // memory_array[25155] <= 3'b111;
      // memory_array[25156] <= 3'b111;
      // memory_array[25157] <= 3'b111;
      // memory_array[25158] <= 3'b111;
      // memory_array[25159] <= 3'b111;
      // memory_array[25160] <= 3'b111;
      // memory_array[25161] <= 3'b000;
      // memory_array[25162] <= 3'b111;
      // memory_array[25163] <= 3'b110;
      // memory_array[25164] <= 3'b110;
      // memory_array[25165] <= 3'b111;
      // memory_array[25166] <= 3'b110;
      // memory_array[25167] <= 3'b111;
      // memory_array[25168] <= 3'b110;
      // memory_array[25169] <= 3'b110;
      // memory_array[25170] <= 3'b110;
      // memory_array[25171] <= 3'b110;
      // memory_array[25172] <= 3'b000;
      // memory_array[25173] <= 3'b110;
      // memory_array[25174] <= 3'b000;
      // memory_array[25175] <= 3'b000;
      // memory_array[25176] <= 3'b111;
      // memory_array[25177] <= 3'b111;
      // memory_array[25178] <= 3'b111;
      // memory_array[25179] <= 3'b000;
      // memory_array[25180] <= 3'b110;
      // memory_array[25181] <= 3'b110;
      // memory_array[25182] <= 3'b110;
      // memory_array[25183] <= 3'b110;
      // memory_array[25184] <= 3'b110;
      // memory_array[25185] <= 3'b000;
      // memory_array[25186] <= 3'b000;
      // memory_array[25187] <= 3'b000;
      // memory_array[25188] <= 3'b110;
      // memory_array[25189] <= 3'b000;
      // memory_array[25190] <= 3'b000;
      // memory_array[25191] <= 3'b101;
      // memory_array[25192] <= 3'b111;
      // memory_array[25193] <= 3'b101;
      // memory_array[25194] <= 3'b101;
      // memory_array[25195] <= 3'b101;
      // memory_array[25196] <= 3'b101;
      // memory_array[25197] <= 3'b101;
      // memory_array[25198] <= 3'b101;
      // memory_array[25199] <= 3'b101;
      // memory_array[25200] <= 3'b101;
      // memory_array[25201] <= 3'b101;
      // memory_array[25202] <= 3'b101;
      // memory_array[25203] <= 3'b111;
      // memory_array[25204] <= 3'b111;
      // memory_array[25205] <= 3'b101;
      // memory_array[25206] <= 3'b101;
      // memory_array[25207] <= 3'b101;
      // memory_array[25208] <= 3'b101;
      // memory_array[25209] <= 3'b000;
      // memory_array[25210] <= 3'b000;
      // memory_array[25211] <= 3'b110;
      // memory_array[25212] <= 3'b000;
      // memory_array[25213] <= 3'b110;
      // memory_array[25214] <= 3'b110;
      // memory_array[25215] <= 3'b000;
      // memory_array[25216] <= 3'b110;
      // memory_array[25217] <= 3'b111;
      // memory_array[25218] <= 3'b110;
      // memory_array[25219] <= 3'b110;
      // memory_array[25220] <= 3'b111;
      // memory_array[25221] <= 3'b000;
      // memory_array[25222] <= 3'b111;
      // memory_array[25223] <= 3'b111;
      // memory_array[25224] <= 3'b000;
      // memory_array[25225] <= 3'b000;
      // memory_array[25226] <= 3'b000;
      // memory_array[25227] <= 3'b110;
      // memory_array[25228] <= 3'b110;
      // memory_array[25229] <= 3'b110;
      // memory_array[25230] <= 3'b111;
      // memory_array[25231] <= 3'b111;
      // memory_array[25232] <= 3'b000;
      // memory_array[25233] <= 3'b110;
      // memory_array[25234] <= 3'b110;
      // memory_array[25235] <= 3'b110;
      // memory_array[25236] <= 3'b110;
      // memory_array[25237] <= 3'b000;
      // memory_array[25238] <= 3'b000;
      // memory_array[25239] <= 3'b111;
      // memory_array[25240] <= 3'b111;
      // memory_array[25241] <= 3'b111;
      // memory_array[25242] <= 3'b111;
      // memory_array[25243] <= 3'b111;
      // memory_array[25244] <= 3'b111;
      // memory_array[25245] <= 3'b111;
      // memory_array[25246] <= 3'b111;
      // memory_array[25247] <= 3'b111;
      // memory_array[25248] <= 3'b111;
      // memory_array[25249] <= 3'b111;
      // memory_array[25250] <= 3'b111;
      // memory_array[25251] <= 3'b111;
      // memory_array[25252] <= 3'b111;
      // memory_array[25253] <= 3'b111;
      // memory_array[25254] <= 3'b101;
      // memory_array[25255] <= 3'b000;
      // memory_array[25256] <= 3'b000;
      // memory_array[25257] <= 3'b000;
      // memory_array[25258] <= 3'b000;
      // memory_array[25259] <= 3'b000;
      // memory_array[25260] <= 3'b000;
      // memory_array[25261] <= 3'b000;
      // memory_array[25262] <= 3'b000;
      // memory_array[25263] <= 3'b000;
      // memory_array[25264] <= 3'b000;
      // memory_array[25265] <= 3'b000;
      // memory_array[25266] <= 3'b000;
      // memory_array[25267] <= 3'b000;
      // memory_array[25268] <= 3'b101;
      // memory_array[25269] <= 3'b101;
      // memory_array[25270] <= 3'b000;
      // memory_array[25271] <= 3'b000;
      // memory_array[25272] <= 3'b000;
      // memory_array[25273] <= 3'b000;
      // memory_array[25274] <= 3'b000;
      // memory_array[25275] <= 3'b000;
      // memory_array[25276] <= 3'b000;
      // memory_array[25277] <= 3'b000;
      // memory_array[25278] <= 3'b101;
      // memory_array[25279] <= 3'b101;
      // memory_array[25280] <= 3'b101;
      // memory_array[25281] <= 3'b000;
      // memory_array[25282] <= 3'b000;
      // memory_array[25283] <= 3'b101;
      // memory_array[25284] <= 3'b101;
      // memory_array[25285] <= 3'b000;
      // memory_array[25286] <= 3'b000;
      // memory_array[25287] <= 3'b000;
      // memory_array[25288] <= 3'b000;
      // memory_array[25289] <= 3'b110;
      // memory_array[25290] <= 3'b000;
      // memory_array[25291] <= 3'b000;
      // memory_array[25292] <= 3'b000;
      // memory_array[25293] <= 3'b110;
      // memory_array[25294] <= 3'b101;
      // memory_array[25295] <= 3'b000;
      // memory_array[25296] <= 3'b000;
      // memory_array[25297] <= 3'b000;
      // memory_array[25298] <= 3'b101;
      // memory_array[25299] <= 3'b000;
      // memory_array[25300] <= 3'b000;
      // memory_array[25301] <= 3'b000;
      // memory_array[25302] <= 3'b000;
      // memory_array[25303] <= 3'b101;
      // memory_array[25304] <= 3'b101;
      // memory_array[25305] <= 3'b000;
      // memory_array[25306] <= 3'b000;
      // memory_array[25307] <= 3'b000;
      // memory_array[25308] <= 3'b000;
      // memory_array[25309] <= 3'b000;
      // memory_array[25310] <= 3'b000;
      // memory_array[25311] <= 3'b000;
      // memory_array[25312] <= 3'b000;
      // memory_array[25313] <= 3'b000;
      // memory_array[25314] <= 3'b101;
      // memory_array[25315] <= 3'b000;
      // memory_array[25316] <= 3'b101;
      // memory_array[25317] <= 3'b000;
      // memory_array[25318] <= 3'b000;
      // memory_array[25319] <= 3'b101;
      // memory_array[25320] <= 3'b000;
      // memory_array[25321] <= 3'b000;
      // memory_array[25322] <= 3'b000;
      // memory_array[25323] <= 3'b000;
      // memory_array[25324] <= 3'b000;
      // memory_array[25325] <= 3'b000;
      // memory_array[25326] <= 3'b000;
      // memory_array[25327] <= 3'b101;
      // memory_array[25328] <= 3'b101;
      // memory_array[25329] <= 3'b000;
      // memory_array[25330] <= 3'b000;
      // memory_array[25331] <= 3'b000;
      // memory_array[25332] <= 3'b000;
      // memory_array[25333] <= 3'b101;
      // memory_array[25334] <= 3'b101;
      // memory_array[25335] <= 3'b000;
      // memory_array[25336] <= 3'b000;
      // memory_array[25337] <= 3'b000;
      // memory_array[25338] <= 3'b000;
      // memory_array[25339] <= 3'b000;
      // memory_array[25340] <= 3'b000;
      // memory_array[25341] <= 3'b000;
      // memory_array[25342] <= 3'b000;
      // memory_array[25343] <= 3'b000;
      // memory_array[25344] <= 3'b000;
      // memory_array[25345] <= 3'b111;
      // memory_array[25346] <= 3'b111;
      // memory_array[25347] <= 3'b111;
      // memory_array[25348] <= 3'b111;
      // memory_array[25349] <= 3'b111;
      // memory_array[25350] <= 3'b111;
      // memory_array[25351] <= 3'b111;
      // memory_array[25352] <= 3'b111;
      // memory_array[25353] <= 3'b111;
      // memory_array[25354] <= 3'b111;
      // memory_array[25355] <= 3'b111;
      // memory_array[25356] <= 3'b111;
      // memory_array[25357] <= 3'b111;
      // memory_array[25358] <= 3'b111;
      // memory_array[25359] <= 3'b111;
      // memory_array[25360] <= 3'b111;
      // memory_array[25361] <= 3'b000;
      // memory_array[25362] <= 3'b111;
      // memory_array[25363] <= 3'b110;
      // memory_array[25364] <= 3'b110;
      // memory_array[25365] <= 3'b111;
      // memory_array[25366] <= 3'b110;
      // memory_array[25367] <= 3'b111;
      // memory_array[25368] <= 3'b110;
      // memory_array[25369] <= 3'b110;
      // memory_array[25370] <= 3'b110;
      // memory_array[25371] <= 3'b110;
      // memory_array[25372] <= 3'b000;
      // memory_array[25373] <= 3'b110;
      // memory_array[25374] <= 3'b110;
      // memory_array[25375] <= 3'b111;
      // memory_array[25376] <= 3'b111;
      // memory_array[25377] <= 3'b000;
      // memory_array[25378] <= 3'b000;
      // memory_array[25379] <= 3'b111;
      // memory_array[25380] <= 3'b111;
      // memory_array[25381] <= 3'b110;
      // memory_array[25382] <= 3'b110;
      // memory_array[25383] <= 3'b110;
      // memory_array[25384] <= 3'b110;
      // memory_array[25385] <= 3'b000;
      // memory_array[25386] <= 3'b000;
      // memory_array[25387] <= 3'b000;
      // memory_array[25388] <= 3'b110;
      // memory_array[25389] <= 3'b000;
      // memory_array[25390] <= 3'b000;
      // memory_array[25391] <= 3'b101;
      // memory_array[25392] <= 3'b101;
      // memory_array[25393] <= 3'b101;
      // memory_array[25394] <= 3'b101;
      // memory_array[25395] <= 3'b111;
      // memory_array[25396] <= 3'b111;
      // memory_array[25397] <= 3'b101;
      // memory_array[25398] <= 3'b101;
      // memory_array[25399] <= 3'b101;
      // memory_array[25400] <= 3'b101;
      // memory_array[25401] <= 3'b000;
      // memory_array[25402] <= 3'b000;
      // memory_array[25403] <= 3'b110;
      // memory_array[25404] <= 3'b110;
      // memory_array[25405] <= 3'b000;
      // memory_array[25406] <= 3'b000;
      // memory_array[25407] <= 3'b101;
      // memory_array[25408] <= 3'b101;
      // memory_array[25409] <= 3'b000;
      // memory_array[25410] <= 3'b000;
      // memory_array[25411] <= 3'b000;
      // memory_array[25412] <= 3'b000;
      // memory_array[25413] <= 3'b000;
      // memory_array[25414] <= 3'b000;
      // memory_array[25415] <= 3'b000;
      // memory_array[25416] <= 3'b000;
      // memory_array[25417] <= 3'b000;
      // memory_array[25418] <= 3'b000;
      // memory_array[25419] <= 3'b000;
      // memory_array[25420] <= 3'b111;
      // memory_array[25421] <= 3'b111;
      // memory_array[25422] <= 3'b000;
      // memory_array[25423] <= 3'b000;
      // memory_array[25424] <= 3'b000;
      // memory_array[25425] <= 3'b000;
      // memory_array[25426] <= 3'b000;
      // memory_array[25427] <= 3'b000;
      // memory_array[25428] <= 3'b000;
      // memory_array[25429] <= 3'b000;
      // memory_array[25430] <= 3'b000;
      // memory_array[25431] <= 3'b000;
      // memory_array[25432] <= 3'b000;
      // memory_array[25433] <= 3'b000;
      // memory_array[25434] <= 3'b000;
      // memory_array[25435] <= 3'b000;
      // memory_array[25436] <= 3'b000;
      // memory_array[25437] <= 3'b000;
      // memory_array[25438] <= 3'b000;
      // memory_array[25439] <= 3'b111;
      // memory_array[25440] <= 3'b111;
      // memory_array[25441] <= 3'b111;
      // memory_array[25442] <= 3'b111;
      // memory_array[25443] <= 3'b111;
      // memory_array[25444] <= 3'b111;
      // memory_array[25445] <= 3'b111;
      // memory_array[25446] <= 3'b111;
      // memory_array[25447] <= 3'b111;
      // memory_array[25448] <= 3'b111;
      // memory_array[25449] <= 3'b111;
      // memory_array[25450] <= 3'b111;
      // memory_array[25451] <= 3'b111;
      // memory_array[25452] <= 3'b111;
      // memory_array[25453] <= 3'b111;
      // memory_array[25454] <= 3'b101;
      // memory_array[25455] <= 3'b000;
      // memory_array[25456] <= 3'b000;
      // memory_array[25457] <= 3'b000;
      // memory_array[25458] <= 3'b000;
      // memory_array[25459] <= 3'b000;
      // memory_array[25460] <= 3'b000;
      // memory_array[25461] <= 3'b000;
      // memory_array[25462] <= 3'b000;
      // memory_array[25463] <= 3'b000;
      // memory_array[25464] <= 3'b000;
      // memory_array[25465] <= 3'b000;
      // memory_array[25466] <= 3'b000;
      // memory_array[25467] <= 3'b000;
      // memory_array[25468] <= 3'b000;
      // memory_array[25469] <= 3'b101;
      // memory_array[25470] <= 3'b000;
      // memory_array[25471] <= 3'b000;
      // memory_array[25472] <= 3'b000;
      // memory_array[25473] <= 3'b101;
      // memory_array[25474] <= 3'b101;
      // memory_array[25475] <= 3'b000;
      // memory_array[25476] <= 3'b000;
      // memory_array[25477] <= 3'b000;
      // memory_array[25478] <= 3'b101;
      // memory_array[25479] <= 3'b000;
      // memory_array[25480] <= 3'b000;
      // memory_array[25481] <= 3'b000;
      // memory_array[25482] <= 3'b000;
      // memory_array[25483] <= 3'b000;
      // memory_array[25484] <= 3'b101;
      // memory_array[25485] <= 3'b000;
      // memory_array[25486] <= 3'b000;
      // memory_array[25487] <= 3'b000;
      // memory_array[25488] <= 3'b000;
      // memory_array[25489] <= 3'b101;
      // memory_array[25490] <= 3'b000;
      // memory_array[25491] <= 3'b000;
      // memory_array[25492] <= 3'b000;
      // memory_array[25493] <= 3'b000;
      // memory_array[25494] <= 3'b110;
      // memory_array[25495] <= 3'b000;
      // memory_array[25496] <= 3'b000;
      // memory_array[25497] <= 3'b000;
      // memory_array[25498] <= 3'b101;
      // memory_array[25499] <= 3'b101;
      // memory_array[25500] <= 3'b000;
      // memory_array[25501] <= 3'b000;
      // memory_array[25502] <= 3'b000;
      // memory_array[25503] <= 3'b000;
      // memory_array[25504] <= 3'b101;
      // memory_array[25505] <= 3'b000;
      // memory_array[25506] <= 3'b000;
      // memory_array[25507] <= 3'b000;
      // memory_array[25508] <= 3'b000;
      // memory_array[25509] <= 3'b000;
      // memory_array[25510] <= 3'b101;
      // memory_array[25511] <= 3'b000;
      // memory_array[25512] <= 3'b000;
      // memory_array[25513] <= 3'b000;
      // memory_array[25514] <= 3'b000;
      // memory_array[25515] <= 3'b000;
      // memory_array[25516] <= 3'b000;
      // memory_array[25517] <= 3'b000;
      // memory_array[25518] <= 3'b000;
      // memory_array[25519] <= 3'b000;
      // memory_array[25520] <= 3'b000;
      // memory_array[25521] <= 3'b000;
      // memory_array[25522] <= 3'b000;
      // memory_array[25523] <= 3'b000;
      // memory_array[25524] <= 3'b000;
      // memory_array[25525] <= 3'b000;
      // memory_array[25526] <= 3'b000;
      // memory_array[25527] <= 3'b000;
      // memory_array[25528] <= 3'b101;
      // memory_array[25529] <= 3'b000;
      // memory_array[25530] <= 3'b000;
      // memory_array[25531] <= 3'b000;
      // memory_array[25532] <= 3'b000;
      // memory_array[25533] <= 3'b101;
      // memory_array[25534] <= 3'b101;
      // memory_array[25535] <= 3'b000;
      // memory_array[25536] <= 3'b000;
      // memory_array[25537] <= 3'b000;
      // memory_array[25538] <= 3'b000;
      // memory_array[25539] <= 3'b000;
      // memory_array[25540] <= 3'b000;
      // memory_array[25541] <= 3'b000;
      // memory_array[25542] <= 3'b000;
      // memory_array[25543] <= 3'b000;
      // memory_array[25544] <= 3'b000;
      // memory_array[25545] <= 3'b111;
      // memory_array[25546] <= 3'b111;
      // memory_array[25547] <= 3'b111;
      // memory_array[25548] <= 3'b111;
      // memory_array[25549] <= 3'b111;
      // memory_array[25550] <= 3'b111;
      // memory_array[25551] <= 3'b111;
      // memory_array[25552] <= 3'b111;
      // memory_array[25553] <= 3'b111;
      // memory_array[25554] <= 3'b111;
      // memory_array[25555] <= 3'b111;
      // memory_array[25556] <= 3'b111;
      // memory_array[25557] <= 3'b111;
      // memory_array[25558] <= 3'b111;
      // memory_array[25559] <= 3'b111;
      // memory_array[25560] <= 3'b111;
      // memory_array[25561] <= 3'b000;
      // memory_array[25562] <= 3'b000;
      // memory_array[25563] <= 3'b000;
      // memory_array[25564] <= 3'b000;
      // memory_array[25565] <= 3'b000;
      // memory_array[25566] <= 3'b000;
      // memory_array[25567] <= 3'b000;
      // memory_array[25568] <= 3'b000;
      // memory_array[25569] <= 3'b000;
      // memory_array[25570] <= 3'b000;
      // memory_array[25571] <= 3'b000;
      // memory_array[25572] <= 3'b000;
      // memory_array[25573] <= 3'b000;
      // memory_array[25574] <= 3'b000;
      // memory_array[25575] <= 3'b000;
      // memory_array[25576] <= 3'b000;
      // memory_array[25577] <= 3'b000;
      // memory_array[25578] <= 3'b000;
      // memory_array[25579] <= 3'b000;
      // memory_array[25580] <= 3'b000;
      // memory_array[25581] <= 3'b111;
      // memory_array[25582] <= 3'b000;
      // memory_array[25583] <= 3'b000;
      // memory_array[25584] <= 3'b000;
      // memory_array[25585] <= 3'b000;
      // memory_array[25586] <= 3'b000;
      // memory_array[25587] <= 3'b000;
      // memory_array[25588] <= 3'b000;
      // memory_array[25589] <= 3'b000;
      // memory_array[25590] <= 3'b000;
      // memory_array[25591] <= 3'b101;
      // memory_array[25592] <= 3'b101;
      // memory_array[25593] <= 3'b110;
      // memory_array[25594] <= 3'b110;
      // memory_array[25595] <= 3'b000;
      // memory_array[25596] <= 3'b000;
      // memory_array[25597] <= 3'b000;
      // memory_array[25598] <= 3'b110;
      // memory_array[25599] <= 3'b101;
      // memory_array[25600] <= 3'b101;
      // memory_array[25601] <= 3'b110;
      // memory_array[25602] <= 3'b110;
      // memory_array[25603] <= 3'b000;
      // memory_array[25604] <= 3'b000;
      // memory_array[25605] <= 3'b110;
      // memory_array[25606] <= 3'b110;
      // memory_array[25607] <= 3'b101;
      // memory_array[25608] <= 3'b101;
      // memory_array[25609] <= 3'b000;
      // memory_array[25610] <= 3'b000;
      // memory_array[25611] <= 3'b000;
      // memory_array[25612] <= 3'b000;
      // memory_array[25613] <= 3'b000;
      // memory_array[25614] <= 3'b000;
      // memory_array[25615] <= 3'b000;
      // memory_array[25616] <= 3'b000;
      // memory_array[25617] <= 3'b000;
      // memory_array[25618] <= 3'b000;
      // memory_array[25619] <= 3'b000;
      // memory_array[25620] <= 3'b000;
      // memory_array[25621] <= 3'b000;
      // memory_array[25622] <= 3'b000;
      // memory_array[25623] <= 3'b000;
      // memory_array[25624] <= 3'b000;
      // memory_array[25625] <= 3'b000;
      // memory_array[25626] <= 3'b000;
      // memory_array[25627] <= 3'b000;
      // memory_array[25628] <= 3'b000;
      // memory_array[25629] <= 3'b000;
      // memory_array[25630] <= 3'b000;
      // memory_array[25631] <= 3'b000;
      // memory_array[25632] <= 3'b000;
      // memory_array[25633] <= 3'b000;
      // memory_array[25634] <= 3'b000;
      // memory_array[25635] <= 3'b000;
      // memory_array[25636] <= 3'b000;
      // memory_array[25637] <= 3'b000;
      // memory_array[25638] <= 3'b000;
      // memory_array[25639] <= 3'b111;
      // memory_array[25640] <= 3'b111;
      // memory_array[25641] <= 3'b111;
      // memory_array[25642] <= 3'b111;
      // memory_array[25643] <= 3'b111;
      // memory_array[25644] <= 3'b111;
      // memory_array[25645] <= 3'b111;
      // memory_array[25646] <= 3'b111;
      // memory_array[25647] <= 3'b111;
      // memory_array[25648] <= 3'b111;
      // memory_array[25649] <= 3'b111;
      // memory_array[25650] <= 3'b111;
      // memory_array[25651] <= 3'b111;
      // memory_array[25652] <= 3'b111;
      // memory_array[25653] <= 3'b111;
      // memory_array[25654] <= 3'b101;
      // memory_array[25655] <= 3'b000;
      // memory_array[25656] <= 3'b000;
      // memory_array[25657] <= 3'b000;
      // memory_array[25658] <= 3'b000;
      // memory_array[25659] <= 3'b000;
      // memory_array[25660] <= 3'b000;
      // memory_array[25661] <= 3'b000;
      // memory_array[25662] <= 3'b000;
      // memory_array[25663] <= 3'b000;
      // memory_array[25664] <= 3'b000;
      // memory_array[25665] <= 3'b000;
      // memory_array[25666] <= 3'b000;
      // memory_array[25667] <= 3'b000;
      // memory_array[25668] <= 3'b000;
      // memory_array[25669] <= 3'b000;
      // memory_array[25670] <= 3'b000;
      // memory_array[25671] <= 3'b000;
      // memory_array[25672] <= 3'b000;
      // memory_array[25673] <= 3'b000;
      // memory_array[25674] <= 3'b000;
      // memory_array[25675] <= 3'b000;
      // memory_array[25676] <= 3'b000;
      // memory_array[25677] <= 3'b000;
      // memory_array[25678] <= 3'b000;
      // memory_array[25679] <= 3'b000;
      // memory_array[25680] <= 3'b000;
      // memory_array[25681] <= 3'b000;
      // memory_array[25682] <= 3'b000;
      // memory_array[25683] <= 3'b000;
      // memory_array[25684] <= 3'b000;
      // memory_array[25685] <= 3'b000;
      // memory_array[25686] <= 3'b000;
      // memory_array[25687] <= 3'b000;
      // memory_array[25688] <= 3'b000;
      // memory_array[25689] <= 3'b000;
      // memory_array[25690] <= 3'b000;
      // memory_array[25691] <= 3'b000;
      // memory_array[25692] <= 3'b000;
      // memory_array[25693] <= 3'b000;
      // memory_array[25694] <= 3'b000;
      // memory_array[25695] <= 3'b000;
      // memory_array[25696] <= 3'b000;
      // memory_array[25697] <= 3'b000;
      // memory_array[25698] <= 3'b000;
      // memory_array[25699] <= 3'b000;
      // memory_array[25700] <= 3'b000;
      // memory_array[25701] <= 3'b000;
      // memory_array[25702] <= 3'b000;
      // memory_array[25703] <= 3'b000;
      // memory_array[25704] <= 3'b000;
      // memory_array[25705] <= 3'b000;
      // memory_array[25706] <= 3'b000;
      // memory_array[25707] <= 3'b000;
      // memory_array[25708] <= 3'b000;
      // memory_array[25709] <= 3'b000;
      // memory_array[25710] <= 3'b000;
      // memory_array[25711] <= 3'b000;
      // memory_array[25712] <= 3'b000;
      // memory_array[25713] <= 3'b000;
      // memory_array[25714] <= 3'b000;
      // memory_array[25715] <= 3'b000;
      // memory_array[25716] <= 3'b000;
      // memory_array[25717] <= 3'b000;
      // memory_array[25718] <= 3'b000;
      // memory_array[25719] <= 3'b000;
      // memory_array[25720] <= 3'b000;
      // memory_array[25721] <= 3'b000;
      // memory_array[25722] <= 3'b000;
      // memory_array[25723] <= 3'b000;
      // memory_array[25724] <= 3'b000;
      // memory_array[25725] <= 3'b000;
      // memory_array[25726] <= 3'b000;
      // memory_array[25727] <= 3'b000;
      // memory_array[25728] <= 3'b000;
      // memory_array[25729] <= 3'b000;
      // memory_array[25730] <= 3'b000;
      // memory_array[25731] <= 3'b000;
      // memory_array[25732] <= 3'b000;
      // memory_array[25733] <= 3'b000;
      // memory_array[25734] <= 3'b000;
      // memory_array[25735] <= 3'b000;
      // memory_array[25736] <= 3'b000;
      // memory_array[25737] <= 3'b000;
      // memory_array[25738] <= 3'b000;
      // memory_array[25739] <= 3'b000;
      // memory_array[25740] <= 3'b000;
      // memory_array[25741] <= 3'b000;
      // memory_array[25742] <= 3'b000;
      // memory_array[25743] <= 3'b000;
      // memory_array[25744] <= 3'b000;
      // memory_array[25745] <= 3'b111;
      // memory_array[25746] <= 3'b111;
      // memory_array[25747] <= 3'b111;
      // memory_array[25748] <= 3'b111;
      // memory_array[25749] <= 3'b111;
      // memory_array[25750] <= 3'b111;
      // memory_array[25751] <= 3'b111;
      // memory_array[25752] <= 3'b111;
      // memory_array[25753] <= 3'b111;
      // memory_array[25754] <= 3'b111;
      // memory_array[25755] <= 3'b111;
      // memory_array[25756] <= 3'b111;
      // memory_array[25757] <= 3'b111;
      // memory_array[25758] <= 3'b111;
      // memory_array[25759] <= 3'b111;
      // memory_array[25760] <= 3'b111;
      // memory_array[25761] <= 3'b000;
      // memory_array[25762] <= 3'b000;
      // memory_array[25763] <= 3'b000;
      // memory_array[25764] <= 3'b000;
      // memory_array[25765] <= 3'b000;
      // memory_array[25766] <= 3'b000;
      // memory_array[25767] <= 3'b000;
      // memory_array[25768] <= 3'b000;
      // memory_array[25769] <= 3'b000;
      // memory_array[25770] <= 3'b000;
      // memory_array[25771] <= 3'b000;
      // memory_array[25772] <= 3'b000;
      // memory_array[25773] <= 3'b000;
      // memory_array[25774] <= 3'b000;
      // memory_array[25775] <= 3'b000;
      // memory_array[25776] <= 3'b000;
      // memory_array[25777] <= 3'b000;
      // memory_array[25778] <= 3'b000;
      // memory_array[25779] <= 3'b000;
      // memory_array[25780] <= 3'b000;
      // memory_array[25781] <= 3'b000;
      // memory_array[25782] <= 3'b000;
      // memory_array[25783] <= 3'b000;
      // memory_array[25784] <= 3'b000;
      // memory_array[25785] <= 3'b000;
      // memory_array[25786] <= 3'b000;
      // memory_array[25787] <= 3'b000;
      // memory_array[25788] <= 3'b000;
      // memory_array[25789] <= 3'b000;
      // memory_array[25790] <= 3'b000;
      // memory_array[25791] <= 3'b101;
      // memory_array[25792] <= 3'b110;
      // memory_array[25793] <= 3'b000;
      // memory_array[25794] <= 3'b000;
      // memory_array[25795] <= 3'b110;
      // memory_array[25796] <= 3'b110;
      // memory_array[25797] <= 3'b110;
      // memory_array[25798] <= 3'b000;
      // memory_array[25799] <= 3'b101;
      // memory_array[25800] <= 3'b000;
      // memory_array[25801] <= 3'b000;
      // memory_array[25802] <= 3'b000;
      // memory_array[25803] <= 3'b110;
      // memory_array[25804] <= 3'b110;
      // memory_array[25805] <= 3'b000;
      // memory_array[25806] <= 3'b000;
      // memory_array[25807] <= 3'b000;
      // memory_array[25808] <= 3'b101;
      // memory_array[25809] <= 3'b000;
      // memory_array[25810] <= 3'b000;
      // memory_array[25811] <= 3'b000;
      // memory_array[25812] <= 3'b000;
      // memory_array[25813] <= 3'b000;
      // memory_array[25814] <= 3'b000;
      // memory_array[25815] <= 3'b000;
      // memory_array[25816] <= 3'b000;
      // memory_array[25817] <= 3'b000;
      // memory_array[25818] <= 3'b000;
      // memory_array[25819] <= 3'b000;
      // memory_array[25820] <= 3'b000;
      // memory_array[25821] <= 3'b000;
      // memory_array[25822] <= 3'b000;
      // memory_array[25823] <= 3'b000;
      // memory_array[25824] <= 3'b000;
      // memory_array[25825] <= 3'b000;
      // memory_array[25826] <= 3'b000;
      // memory_array[25827] <= 3'b000;
      // memory_array[25828] <= 3'b000;
      // memory_array[25829] <= 3'b000;
      // memory_array[25830] <= 3'b000;
      // memory_array[25831] <= 3'b000;
      // memory_array[25832] <= 3'b000;
      // memory_array[25833] <= 3'b000;
      // memory_array[25834] <= 3'b000;
      // memory_array[25835] <= 3'b000;
      // memory_array[25836] <= 3'b000;
      // memory_array[25837] <= 3'b000;
      // memory_array[25838] <= 3'b000;
      // memory_array[25839] <= 3'b111;
      // memory_array[25840] <= 3'b111;
      // memory_array[25841] <= 3'b111;
      // memory_array[25842] <= 3'b111;
      // memory_array[25843] <= 3'b111;
      // memory_array[25844] <= 3'b111;
      // memory_array[25845] <= 3'b111;
      // memory_array[25846] <= 3'b111;
      // memory_array[25847] <= 3'b111;
      // memory_array[25848] <= 3'b111;
      // memory_array[25849] <= 3'b111;
      // memory_array[25850] <= 3'b111;
      // memory_array[25851] <= 3'b111;
      // memory_array[25852] <= 3'b111;
      // memory_array[25853] <= 3'b111;
      // memory_array[25854] <= 3'b101;
      // memory_array[25855] <= 3'b000;
      // memory_array[25856] <= 3'b000;
      // memory_array[25857] <= 3'b000;
      // memory_array[25858] <= 3'b000;
      // memory_array[25859] <= 3'b000;
      // memory_array[25860] <= 3'b000;
      // memory_array[25861] <= 3'b000;
      // memory_array[25862] <= 3'b000;
      // memory_array[25863] <= 3'b000;
      // memory_array[25864] <= 3'b000;
      // memory_array[25865] <= 3'b000;
      // memory_array[25866] <= 3'b000;
      // memory_array[25867] <= 3'b000;
      // memory_array[25868] <= 3'b000;
      // memory_array[25869] <= 3'b000;
      // memory_array[25870] <= 3'b000;
      // memory_array[25871] <= 3'b000;
      // memory_array[25872] <= 3'b000;
      // memory_array[25873] <= 3'b000;
      // memory_array[25874] <= 3'b000;
      // memory_array[25875] <= 3'b000;
      // memory_array[25876] <= 3'b000;
      // memory_array[25877] <= 3'b000;
      // memory_array[25878] <= 3'b000;
      // memory_array[25879] <= 3'b000;
      // memory_array[25880] <= 3'b000;
      // memory_array[25881] <= 3'b000;
      // memory_array[25882] <= 3'b000;
      // memory_array[25883] <= 3'b000;
      // memory_array[25884] <= 3'b000;
      // memory_array[25885] <= 3'b000;
      // memory_array[25886] <= 3'b000;
      // memory_array[25887] <= 3'b000;
      // memory_array[25888] <= 3'b000;
      // memory_array[25889] <= 3'b000;
      // memory_array[25890] <= 3'b000;
      // memory_array[25891] <= 3'b000;
      // memory_array[25892] <= 3'b000;
      // memory_array[25893] <= 3'b000;
      // memory_array[25894] <= 3'b000;
      // memory_array[25895] <= 3'b000;
      // memory_array[25896] <= 3'b000;
      // memory_array[25897] <= 3'b000;
      // memory_array[25898] <= 3'b000;
      // memory_array[25899] <= 3'b000;
      // memory_array[25900] <= 3'b000;
      // memory_array[25901] <= 3'b000;
      // memory_array[25902] <= 3'b000;
      // memory_array[25903] <= 3'b000;
      // memory_array[25904] <= 3'b000;
      // memory_array[25905] <= 3'b000;
      // memory_array[25906] <= 3'b000;
      // memory_array[25907] <= 3'b000;
      // memory_array[25908] <= 3'b000;
      // memory_array[25909] <= 3'b000;
      // memory_array[25910] <= 3'b000;
      // memory_array[25911] <= 3'b000;
      // memory_array[25912] <= 3'b000;
      // memory_array[25913] <= 3'b000;
      // memory_array[25914] <= 3'b000;
      // memory_array[25915] <= 3'b000;
      // memory_array[25916] <= 3'b000;
      // memory_array[25917] <= 3'b000;
      // memory_array[25918] <= 3'b000;
      // memory_array[25919] <= 3'b000;
      // memory_array[25920] <= 3'b000;
      // memory_array[25921] <= 3'b000;
      // memory_array[25922] <= 3'b000;
      // memory_array[25923] <= 3'b000;
      // memory_array[25924] <= 3'b000;
      // memory_array[25925] <= 3'b000;
      // memory_array[25926] <= 3'b000;
      // memory_array[25927] <= 3'b000;
      // memory_array[25928] <= 3'b000;
      // memory_array[25929] <= 3'b000;
      // memory_array[25930] <= 3'b000;
      // memory_array[25931] <= 3'b000;
      // memory_array[25932] <= 3'b000;
      // memory_array[25933] <= 3'b000;
      // memory_array[25934] <= 3'b000;
      // memory_array[25935] <= 3'b000;
      // memory_array[25936] <= 3'b000;
      // memory_array[25937] <= 3'b000;
      // memory_array[25938] <= 3'b000;
      // memory_array[25939] <= 3'b000;
      // memory_array[25940] <= 3'b000;
      // memory_array[25941] <= 3'b000;
      // memory_array[25942] <= 3'b000;
      // memory_array[25943] <= 3'b000;
      // memory_array[25944] <= 3'b000;
      // memory_array[25945] <= 3'b111;
      // memory_array[25946] <= 3'b111;
      // memory_array[25947] <= 3'b111;
      // memory_array[25948] <= 3'b111;
      // memory_array[25949] <= 3'b111;
      // memory_array[25950] <= 3'b111;
      // memory_array[25951] <= 3'b111;
      // memory_array[25952] <= 3'b111;
      // memory_array[25953] <= 3'b111;
      // memory_array[25954] <= 3'b111;
      // memory_array[25955] <= 3'b111;
      // memory_array[25956] <= 3'b111;
      // memory_array[25957] <= 3'b111;
      // memory_array[25958] <= 3'b111;
      // memory_array[25959] <= 3'b111;
      // memory_array[25960] <= 3'b111;
      // memory_array[25961] <= 3'b000;
      // memory_array[25962] <= 3'b000;
      // memory_array[25963] <= 3'b000;
      // memory_array[25964] <= 3'b000;
      // memory_array[25965] <= 3'b000;
      // memory_array[25966] <= 3'b000;
      // memory_array[25967] <= 3'b000;
      // memory_array[25968] <= 3'b000;
      // memory_array[25969] <= 3'b000;
      // memory_array[25970] <= 3'b000;
      // memory_array[25971] <= 3'b000;
      // memory_array[25972] <= 3'b000;
      // memory_array[25973] <= 3'b000;
      // memory_array[25974] <= 3'b000;
      // memory_array[25975] <= 3'b000;
      // memory_array[25976] <= 3'b000;
      // memory_array[25977] <= 3'b000;
      // memory_array[25978] <= 3'b000;
      // memory_array[25979] <= 3'b000;
      // memory_array[25980] <= 3'b000;
      // memory_array[25981] <= 3'b000;
      // memory_array[25982] <= 3'b000;
      // memory_array[25983] <= 3'b000;
      // memory_array[25984] <= 3'b000;
      // memory_array[25985] <= 3'b000;
      // memory_array[25986] <= 3'b000;
      // memory_array[25987] <= 3'b000;
      // memory_array[25988] <= 3'b000;
      // memory_array[25989] <= 3'b000;
      // memory_array[25990] <= 3'b000;
      // memory_array[25991] <= 3'b101;
      // memory_array[25992] <= 3'b000;
      // memory_array[25993] <= 3'b110;
      // memory_array[25994] <= 3'b110;
      // memory_array[25995] <= 3'b000;
      // memory_array[25996] <= 3'b000;
      // memory_array[25997] <= 3'b000;
      // memory_array[25998] <= 3'b110;
      // memory_array[25999] <= 3'b110;
      // memory_array[26000] <= 3'b101;
      // memory_array[26001] <= 3'b101;
      // memory_array[26002] <= 3'b101;
      // memory_array[26003] <= 3'b101;
      // memory_array[26004] <= 3'b101;
      // memory_array[26005] <= 3'b101;
      // memory_array[26006] <= 3'b101;
      // memory_array[26007] <= 3'b101;
      // memory_array[26008] <= 3'b101;
      // memory_array[26009] <= 3'b000;
      // memory_array[26010] <= 3'b000;
      // memory_array[26011] <= 3'b000;
      // memory_array[26012] <= 3'b000;
      // memory_array[26013] <= 3'b000;
      // memory_array[26014] <= 3'b000;
      // memory_array[26015] <= 3'b000;
      // memory_array[26016] <= 3'b000;
      // memory_array[26017] <= 3'b000;
      // memory_array[26018] <= 3'b000;
      // memory_array[26019] <= 3'b000;
      // memory_array[26020] <= 3'b000;
      // memory_array[26021] <= 3'b000;
      // memory_array[26022] <= 3'b000;
      // memory_array[26023] <= 3'b000;
      // memory_array[26024] <= 3'b000;
      // memory_array[26025] <= 3'b000;
      // memory_array[26026] <= 3'b000;
      // memory_array[26027] <= 3'b000;
      // memory_array[26028] <= 3'b000;
      // memory_array[26029] <= 3'b000;
      // memory_array[26030] <= 3'b000;
      // memory_array[26031] <= 3'b000;
      // memory_array[26032] <= 3'b000;
      // memory_array[26033] <= 3'b000;
      // memory_array[26034] <= 3'b000;
      // memory_array[26035] <= 3'b000;
      // memory_array[26036] <= 3'b000;
      // memory_array[26037] <= 3'b000;
      // memory_array[26038] <= 3'b000;
      // memory_array[26039] <= 3'b111;
      // memory_array[26040] <= 3'b111;
      // memory_array[26041] <= 3'b111;
      // memory_array[26042] <= 3'b111;
      // memory_array[26043] <= 3'b111;
      // memory_array[26044] <= 3'b111;
      // memory_array[26045] <= 3'b111;
      // memory_array[26046] <= 3'b111;
      // memory_array[26047] <= 3'b111;
      // memory_array[26048] <= 3'b111;
      // memory_array[26049] <= 3'b111;
      // memory_array[26050] <= 3'b111;
      // memory_array[26051] <= 3'b111;
      // memory_array[26052] <= 3'b111;
      // memory_array[26053] <= 3'b111;
      // memory_array[26054] <= 3'b101;
      // memory_array[26055] <= 3'b000;
      // memory_array[26056] <= 3'b000;
      // memory_array[26057] <= 3'b000;
      // memory_array[26058] <= 3'b000;
      // memory_array[26059] <= 3'b000;
      // memory_array[26060] <= 3'b000;
      // memory_array[26061] <= 3'b000;
      // memory_array[26062] <= 3'b000;
      // memory_array[26063] <= 3'b000;
      // memory_array[26064] <= 3'b000;
      // memory_array[26065] <= 3'b000;
      // memory_array[26066] <= 3'b000;
      // memory_array[26067] <= 3'b000;
      // memory_array[26068] <= 3'b000;
      // memory_array[26069] <= 3'b000;
      // memory_array[26070] <= 3'b000;
      // memory_array[26071] <= 3'b000;
      // memory_array[26072] <= 3'b000;
      // memory_array[26073] <= 3'b000;
      // memory_array[26074] <= 3'b000;
      // memory_array[26075] <= 3'b000;
      // memory_array[26076] <= 3'b000;
      // memory_array[26077] <= 3'b000;
      // memory_array[26078] <= 3'b000;
      // memory_array[26079] <= 3'b000;
      // memory_array[26080] <= 3'b000;
      // memory_array[26081] <= 3'b000;
      // memory_array[26082] <= 3'b000;
      // memory_array[26083] <= 3'b000;
      // memory_array[26084] <= 3'b000;
      // memory_array[26085] <= 3'b000;
      // memory_array[26086] <= 3'b000;
      // memory_array[26087] <= 3'b000;
      // memory_array[26088] <= 3'b000;
      // memory_array[26089] <= 3'b000;
      // memory_array[26090] <= 3'b000;
      // memory_array[26091] <= 3'b000;
      // memory_array[26092] <= 3'b000;
      // memory_array[26093] <= 3'b000;
      // memory_array[26094] <= 3'b000;
      // memory_array[26095] <= 3'b000;
      // memory_array[26096] <= 3'b000;
      // memory_array[26097] <= 3'b000;
      // memory_array[26098] <= 3'b000;
      // memory_array[26099] <= 3'b000;
      // memory_array[26100] <= 3'b000;
      // memory_array[26101] <= 3'b000;
      // memory_array[26102] <= 3'b000;
      // memory_array[26103] <= 3'b000;
      // memory_array[26104] <= 3'b000;
      // memory_array[26105] <= 3'b000;
      // memory_array[26106] <= 3'b000;
      // memory_array[26107] <= 3'b000;
      // memory_array[26108] <= 3'b000;
      // memory_array[26109] <= 3'b000;
      // memory_array[26110] <= 3'b000;
      // memory_array[26111] <= 3'b000;
      // memory_array[26112] <= 3'b000;
      // memory_array[26113] <= 3'b000;
      // memory_array[26114] <= 3'b000;
      // memory_array[26115] <= 3'b000;
      // memory_array[26116] <= 3'b000;
      // memory_array[26117] <= 3'b000;
      // memory_array[26118] <= 3'b000;
      // memory_array[26119] <= 3'b000;
      // memory_array[26120] <= 3'b000;
      // memory_array[26121] <= 3'b000;
      // memory_array[26122] <= 3'b000;
      // memory_array[26123] <= 3'b000;
      // memory_array[26124] <= 3'b000;
      // memory_array[26125] <= 3'b000;
      // memory_array[26126] <= 3'b000;
      // memory_array[26127] <= 3'b000;
      // memory_array[26128] <= 3'b000;
      // memory_array[26129] <= 3'b000;
      // memory_array[26130] <= 3'b000;
      // memory_array[26131] <= 3'b000;
      // memory_array[26132] <= 3'b000;
      // memory_array[26133] <= 3'b000;
      // memory_array[26134] <= 3'b000;
      // memory_array[26135] <= 3'b000;
      // memory_array[26136] <= 3'b000;
      // memory_array[26137] <= 3'b000;
      // memory_array[26138] <= 3'b000;
      // memory_array[26139] <= 3'b000;
      // memory_array[26140] <= 3'b000;
      // memory_array[26141] <= 3'b000;
      // memory_array[26142] <= 3'b000;
      // memory_array[26143] <= 3'b000;
      // memory_array[26144] <= 3'b000;
      // memory_array[26145] <= 3'b111;
      // memory_array[26146] <= 3'b111;
      // memory_array[26147] <= 3'b111;
      // memory_array[26148] <= 3'b111;
      // memory_array[26149] <= 3'b111;
      // memory_array[26150] <= 3'b111;
      // memory_array[26151] <= 3'b111;
      // memory_array[26152] <= 3'b111;
      // memory_array[26153] <= 3'b111;
      // memory_array[26154] <= 3'b111;
      // memory_array[26155] <= 3'b111;
      // memory_array[26156] <= 3'b111;
      // memory_array[26157] <= 3'b111;
      // memory_array[26158] <= 3'b111;
      // memory_array[26159] <= 3'b111;
      // memory_array[26160] <= 3'b111;
      // memory_array[26161] <= 3'b000;
      // memory_array[26162] <= 3'b000;
      // memory_array[26163] <= 3'b000;
      // memory_array[26164] <= 3'b000;
      // memory_array[26165] <= 3'b000;
      // memory_array[26166] <= 3'b000;
      // memory_array[26167] <= 3'b000;
      // memory_array[26168] <= 3'b000;
      // memory_array[26169] <= 3'b000;
      // memory_array[26170] <= 3'b000;
      // memory_array[26171] <= 3'b000;
      // memory_array[26172] <= 3'b000;
      // memory_array[26173] <= 3'b000;
      // memory_array[26174] <= 3'b000;
      // memory_array[26175] <= 3'b000;
      // memory_array[26176] <= 3'b000;
      // memory_array[26177] <= 3'b000;
      // memory_array[26178] <= 3'b000;
      // memory_array[26179] <= 3'b000;
      // memory_array[26180] <= 3'b000;
      // memory_array[26181] <= 3'b000;
      // memory_array[26182] <= 3'b000;
      // memory_array[26183] <= 3'b000;
      // memory_array[26184] <= 3'b000;
      // memory_array[26185] <= 3'b000;
      // memory_array[26186] <= 3'b000;
      // memory_array[26187] <= 3'b000;
      // memory_array[26188] <= 3'b000;
      // memory_array[26189] <= 3'b000;
      // memory_array[26190] <= 3'b000;
      // memory_array[26191] <= 3'b101;
      // memory_array[26192] <= 3'b101;
      // memory_array[26193] <= 3'b101;
      // memory_array[26194] <= 3'b101;
      // memory_array[26195] <= 3'b101;
      // memory_array[26196] <= 3'b101;
      // memory_array[26197] <= 3'b101;
      // memory_array[26198] <= 3'b101;
      // memory_array[26199] <= 3'b101;
      // memory_array[26200] <= 3'b101;
      // memory_array[26201] <= 3'b101;
      // memory_array[26202] <= 3'b101;
      // memory_array[26203] <= 3'b101;
      // memory_array[26204] <= 3'b101;
      // memory_array[26205] <= 3'b101;
      // memory_array[26206] <= 3'b101;
      // memory_array[26207] <= 3'b101;
      // memory_array[26208] <= 3'b101;
      // memory_array[26209] <= 3'b111;
      // memory_array[26210] <= 3'b111;
      // memory_array[26211] <= 3'b111;
      // memory_array[26212] <= 3'b111;
      // memory_array[26213] <= 3'b111;
      // memory_array[26214] <= 3'b111;
      // memory_array[26215] <= 3'b111;
      // memory_array[26216] <= 3'b111;
      // memory_array[26217] <= 3'b111;
      // memory_array[26218] <= 3'b111;
      // memory_array[26219] <= 3'b111;
      // memory_array[26220] <= 3'b111;
      // memory_array[26221] <= 3'b111;
      // memory_array[26222] <= 3'b111;
      // memory_array[26223] <= 3'b111;
      // memory_array[26224] <= 3'b111;
      // memory_array[26225] <= 3'b111;
      // memory_array[26226] <= 3'b111;
      // memory_array[26227] <= 3'b111;
      // memory_array[26228] <= 3'b111;
      // memory_array[26229] <= 3'b111;
      // memory_array[26230] <= 3'b111;
      // memory_array[26231] <= 3'b111;
      // memory_array[26232] <= 3'b111;
      // memory_array[26233] <= 3'b111;
      // memory_array[26234] <= 3'b111;
      // memory_array[26235] <= 3'b111;
      // memory_array[26236] <= 3'b111;
      // memory_array[26237] <= 3'b111;
      // memory_array[26238] <= 3'b101;
      // memory_array[26239] <= 3'b111;
      // memory_array[26240] <= 3'b111;
      // memory_array[26241] <= 3'b111;
      // memory_array[26242] <= 3'b111;
      // memory_array[26243] <= 3'b111;
      // memory_array[26244] <= 3'b111;
      // memory_array[26245] <= 3'b111;
      // memory_array[26246] <= 3'b111;
      // memory_array[26247] <= 3'b111;
      // memory_array[26248] <= 3'b111;
      // memory_array[26249] <= 3'b111;
      // memory_array[26250] <= 3'b111;
      // memory_array[26251] <= 3'b111;
      // memory_array[26252] <= 3'b111;
      // memory_array[26253] <= 3'b111;
      // memory_array[26254] <= 3'b101;
      // memory_array[26255] <= 3'b101;
      // memory_array[26256] <= 3'b111;
      // memory_array[26257] <= 3'b111;
      // memory_array[26258] <= 3'b111;
      // memory_array[26259] <= 3'b111;
      // memory_array[26260] <= 3'b111;
      // memory_array[26261] <= 3'b111;
      // memory_array[26262] <= 3'b111;
      // memory_array[26263] <= 3'b111;
      // memory_array[26264] <= 3'b111;
      // memory_array[26265] <= 3'b111;
      // memory_array[26266] <= 3'b111;
      // memory_array[26267] <= 3'b111;
      // memory_array[26268] <= 3'b111;
      // memory_array[26269] <= 3'b111;
      // memory_array[26270] <= 3'b111;
      // memory_array[26271] <= 3'b111;
      // memory_array[26272] <= 3'b111;
      // memory_array[26273] <= 3'b111;
      // memory_array[26274] <= 3'b111;
      // memory_array[26275] <= 3'b111;
      // memory_array[26276] <= 3'b111;
      // memory_array[26277] <= 3'b111;
      // memory_array[26278] <= 3'b111;
      // memory_array[26279] <= 3'b111;
      // memory_array[26280] <= 3'b111;
      // memory_array[26281] <= 3'b111;
      // memory_array[26282] <= 3'b111;
      // memory_array[26283] <= 3'b111;
      // memory_array[26284] <= 3'b111;
      // memory_array[26285] <= 3'b111;
      // memory_array[26286] <= 3'b111;
      // memory_array[26287] <= 3'b111;
      // memory_array[26288] <= 3'b111;
      // memory_array[26289] <= 3'b111;
      // memory_array[26290] <= 3'b111;
      // memory_array[26291] <= 3'b111;
      // memory_array[26292] <= 3'b111;
      // memory_array[26293] <= 3'b111;
      // memory_array[26294] <= 3'b111;
      // memory_array[26295] <= 3'b111;
      // memory_array[26296] <= 3'b111;
      // memory_array[26297] <= 3'b111;
      // memory_array[26298] <= 3'b111;
      // memory_array[26299] <= 3'b111;
      // memory_array[26300] <= 3'b111;
      // memory_array[26301] <= 3'b111;
      // memory_array[26302] <= 3'b111;
      // memory_array[26303] <= 3'b111;
      // memory_array[26304] <= 3'b111;
      // memory_array[26305] <= 3'b111;
      // memory_array[26306] <= 3'b111;
      // memory_array[26307] <= 3'b111;
      // memory_array[26308] <= 3'b111;
      // memory_array[26309] <= 3'b111;
      // memory_array[26310] <= 3'b111;
      // memory_array[26311] <= 3'b111;
      // memory_array[26312] <= 3'b111;
      // memory_array[26313] <= 3'b111;
      // memory_array[26314] <= 3'b111;
      // memory_array[26315] <= 3'b111;
      // memory_array[26316] <= 3'b111;
      // memory_array[26317] <= 3'b111;
      // memory_array[26318] <= 3'b111;
      // memory_array[26319] <= 3'b111;
      // memory_array[26320] <= 3'b111;
      // memory_array[26321] <= 3'b111;
      // memory_array[26322] <= 3'b111;
      // memory_array[26323] <= 3'b111;
      // memory_array[26324] <= 3'b111;
      // memory_array[26325] <= 3'b111;
      // memory_array[26326] <= 3'b111;
      // memory_array[26327] <= 3'b111;
      // memory_array[26328] <= 3'b111;
      // memory_array[26329] <= 3'b111;
      // memory_array[26330] <= 3'b111;
      // memory_array[26331] <= 3'b111;
      // memory_array[26332] <= 3'b111;
      // memory_array[26333] <= 3'b111;
      // memory_array[26334] <= 3'b111;
      // memory_array[26335] <= 3'b111;
      // memory_array[26336] <= 3'b111;
      // memory_array[26337] <= 3'b111;
      // memory_array[26338] <= 3'b111;
      // memory_array[26339] <= 3'b111;
      // memory_array[26340] <= 3'b111;
      // memory_array[26341] <= 3'b111;
      // memory_array[26342] <= 3'b111;
      // memory_array[26343] <= 3'b111;
      // memory_array[26344] <= 3'b101;
      // memory_array[26345] <= 3'b111;
      // memory_array[26346] <= 3'b111;
      // memory_array[26347] <= 3'b111;
      // memory_array[26348] <= 3'b111;
      // memory_array[26349] <= 3'b111;
      // memory_array[26350] <= 3'b111;
      // memory_array[26351] <= 3'b111;
      // memory_array[26352] <= 3'b111;
      // memory_array[26353] <= 3'b111;
      // memory_array[26354] <= 3'b111;
      // memory_array[26355] <= 3'b111;
      // memory_array[26356] <= 3'b111;
      // memory_array[26357] <= 3'b111;
      // memory_array[26358] <= 3'b111;
      // memory_array[26359] <= 3'b111;
      // memory_array[26360] <= 3'b111;
      // memory_array[26361] <= 3'b101;
      // memory_array[26362] <= 3'b111;
      // memory_array[26363] <= 3'b111;
      // memory_array[26364] <= 3'b111;
      // memory_array[26365] <= 3'b111;
      // memory_array[26366] <= 3'b111;
      // memory_array[26367] <= 3'b111;
      // memory_array[26368] <= 3'b111;
      // memory_array[26369] <= 3'b111;
      // memory_array[26370] <= 3'b111;
      // memory_array[26371] <= 3'b111;
      // memory_array[26372] <= 3'b111;
      // memory_array[26373] <= 3'b111;
      // memory_array[26374] <= 3'b111;
      // memory_array[26375] <= 3'b111;
      // memory_array[26376] <= 3'b111;
      // memory_array[26377] <= 3'b111;
      // memory_array[26378] <= 3'b111;
      // memory_array[26379] <= 3'b111;
      // memory_array[26380] <= 3'b111;
      // memory_array[26381] <= 3'b111;
      // memory_array[26382] <= 3'b111;
      // memory_array[26383] <= 3'b111;
      // memory_array[26384] <= 3'b111;
      // memory_array[26385] <= 3'b111;
      // memory_array[26386] <= 3'b111;
      // memory_array[26387] <= 3'b111;
      // memory_array[26388] <= 3'b111;
      // memory_array[26389] <= 3'b111;
      // memory_array[26390] <= 3'b111;
      // memory_array[26391] <= 3'b101;
      // memory_array[26392] <= 3'b101;
      // memory_array[26393] <= 3'b101;
      // memory_array[26394] <= 3'b101;
      // memory_array[26395] <= 3'b101;
      // memory_array[26396] <= 3'b101;
      // memory_array[26397] <= 3'b101;
      // memory_array[26398] <= 3'b101;
      // memory_array[26399] <= 3'b101;
      // memory_array[26400] <= 3'b111;
      // memory_array[26401] <= 3'b111;
      // memory_array[26402] <= 3'b111;
      // memory_array[26403] <= 3'b111;
      // memory_array[26404] <= 3'b111;
      // memory_array[26405] <= 3'b111;
      // memory_array[26406] <= 3'b111;
      // memory_array[26407] <= 3'b111;
      // memory_array[26408] <= 3'b101;
      // memory_array[26409] <= 3'b101;
      // memory_array[26410] <= 3'b101;
      // memory_array[26411] <= 3'b101;
      // memory_array[26412] <= 3'b101;
      // memory_array[26413] <= 3'b101;
      // memory_array[26414] <= 3'b101;
      // memory_array[26415] <= 3'b101;
      // memory_array[26416] <= 3'b101;
      // memory_array[26417] <= 3'b101;
      // memory_array[26418] <= 3'b101;
      // memory_array[26419] <= 3'b101;
      // memory_array[26420] <= 3'b101;
      // memory_array[26421] <= 3'b101;
      // memory_array[26422] <= 3'b101;
      // memory_array[26423] <= 3'b101;
      // memory_array[26424] <= 3'b101;
      // memory_array[26425] <= 3'b101;
      // memory_array[26426] <= 3'b101;
      // memory_array[26427] <= 3'b101;
      // memory_array[26428] <= 3'b101;
      // memory_array[26429] <= 3'b101;
      // memory_array[26430] <= 3'b101;
      // memory_array[26431] <= 3'b101;
      // memory_array[26432] <= 3'b101;
      // memory_array[26433] <= 3'b101;
      // memory_array[26434] <= 3'b101;
      // memory_array[26435] <= 3'b101;
      // memory_array[26436] <= 3'b101;
      // memory_array[26437] <= 3'b101;
      // memory_array[26438] <= 3'b101;
      // memory_array[26439] <= 3'b101;
      // memory_array[26440] <= 3'b101;
      // memory_array[26441] <= 3'b101;
      // memory_array[26442] <= 3'b101;
      // memory_array[26443] <= 3'b101;
      // memory_array[26444] <= 3'b101;
      // memory_array[26445] <= 3'b101;
      // memory_array[26446] <= 3'b101;
      // memory_array[26447] <= 3'b101;
      // memory_array[26448] <= 3'b101;
      // memory_array[26449] <= 3'b101;
      // memory_array[26450] <= 3'b101;
      // memory_array[26451] <= 3'b101;
      // memory_array[26452] <= 3'b101;
      // memory_array[26453] <= 3'b101;
      // memory_array[26454] <= 3'b101;
      // memory_array[26455] <= 3'b101;
      // memory_array[26456] <= 3'b101;
      // memory_array[26457] <= 3'b101;
      // memory_array[26458] <= 3'b101;
      // memory_array[26459] <= 3'b101;
      // memory_array[26460] <= 3'b101;
      // memory_array[26461] <= 3'b101;
      // memory_array[26462] <= 3'b101;
      // memory_array[26463] <= 3'b101;
      // memory_array[26464] <= 3'b101;
      // memory_array[26465] <= 3'b101;
      // memory_array[26466] <= 3'b101;
      // memory_array[26467] <= 3'b101;
      // memory_array[26468] <= 3'b101;
      // memory_array[26469] <= 3'b101;
      // memory_array[26470] <= 3'b101;
      // memory_array[26471] <= 3'b101;
      // memory_array[26472] <= 3'b101;
      // memory_array[26473] <= 3'b101;
      // memory_array[26474] <= 3'b101;
      // memory_array[26475] <= 3'b101;
      // memory_array[26476] <= 3'b101;
      // memory_array[26477] <= 3'b101;
      // memory_array[26478] <= 3'b101;
      // memory_array[26479] <= 3'b101;
      // memory_array[26480] <= 3'b101;
      // memory_array[26481] <= 3'b101;
      // memory_array[26482] <= 3'b101;
      // memory_array[26483] <= 3'b101;
      // memory_array[26484] <= 3'b101;
      // memory_array[26485] <= 3'b101;
      // memory_array[26486] <= 3'b101;
      // memory_array[26487] <= 3'b101;
      // memory_array[26488] <= 3'b101;
      // memory_array[26489] <= 3'b101;
      // memory_array[26490] <= 3'b101;
      // memory_array[26491] <= 3'b101;
      // memory_array[26492] <= 3'b101;
      // memory_array[26493] <= 3'b101;
      // memory_array[26494] <= 3'b101;
      // memory_array[26495] <= 3'b101;
      // memory_array[26496] <= 3'b101;
      // memory_array[26497] <= 3'b101;
      // memory_array[26498] <= 3'b101;
      // memory_array[26499] <= 3'b101;
      // memory_array[26500] <= 3'b101;
      // memory_array[26501] <= 3'b101;
      // memory_array[26502] <= 3'b101;
      // memory_array[26503] <= 3'b101;
      // memory_array[26504] <= 3'b101;
      // memory_array[26505] <= 3'b101;
      // memory_array[26506] <= 3'b101;
      // memory_array[26507] <= 3'b101;
      // memory_array[26508] <= 3'b101;
      // memory_array[26509] <= 3'b101;
      // memory_array[26510] <= 3'b101;
      // memory_array[26511] <= 3'b101;
      // memory_array[26512] <= 3'b101;
      // memory_array[26513] <= 3'b101;
      // memory_array[26514] <= 3'b101;
      // memory_array[26515] <= 3'b101;
      // memory_array[26516] <= 3'b101;
      // memory_array[26517] <= 3'b101;
      // memory_array[26518] <= 3'b101;
      // memory_array[26519] <= 3'b101;
      // memory_array[26520] <= 3'b101;
      // memory_array[26521] <= 3'b101;
      // memory_array[26522] <= 3'b101;
      // memory_array[26523] <= 3'b101;
      // memory_array[26524] <= 3'b101;
      // memory_array[26525] <= 3'b101;
      // memory_array[26526] <= 3'b101;
      // memory_array[26527] <= 3'b101;
      // memory_array[26528] <= 3'b101;
      // memory_array[26529] <= 3'b101;
      // memory_array[26530] <= 3'b101;
      // memory_array[26531] <= 3'b101;
      // memory_array[26532] <= 3'b101;
      // memory_array[26533] <= 3'b101;
      // memory_array[26534] <= 3'b101;
      // memory_array[26535] <= 3'b101;
      // memory_array[26536] <= 3'b101;
      // memory_array[26537] <= 3'b101;
      // memory_array[26538] <= 3'b101;
      // memory_array[26539] <= 3'b101;
      // memory_array[26540] <= 3'b101;
      // memory_array[26541] <= 3'b101;
      // memory_array[26542] <= 3'b101;
      // memory_array[26543] <= 3'b101;
      // memory_array[26544] <= 3'b101;
      // memory_array[26545] <= 3'b101;
      // memory_array[26546] <= 3'b101;
      // memory_array[26547] <= 3'b101;
      // memory_array[26548] <= 3'b101;
      // memory_array[26549] <= 3'b101;
      // memory_array[26550] <= 3'b101;
      // memory_array[26551] <= 3'b101;
      // memory_array[26552] <= 3'b101;
      // memory_array[26553] <= 3'b101;
      // memory_array[26554] <= 3'b101;
      // memory_array[26555] <= 3'b101;
      // memory_array[26556] <= 3'b101;
      // memory_array[26557] <= 3'b101;
      // memory_array[26558] <= 3'b101;
      // memory_array[26559] <= 3'b101;
      // memory_array[26560] <= 3'b101;
      // memory_array[26561] <= 3'b101;
      // memory_array[26562] <= 3'b101;
      // memory_array[26563] <= 3'b101;
      // memory_array[26564] <= 3'b101;
      // memory_array[26565] <= 3'b101;
      // memory_array[26566] <= 3'b101;
      // memory_array[26567] <= 3'b101;
      // memory_array[26568] <= 3'b101;
      // memory_array[26569] <= 3'b101;
      // memory_array[26570] <= 3'b101;
      // memory_array[26571] <= 3'b101;
      // memory_array[26572] <= 3'b101;
      // memory_array[26573] <= 3'b101;
      // memory_array[26574] <= 3'b101;
      // memory_array[26575] <= 3'b101;
      // memory_array[26576] <= 3'b101;
      // memory_array[26577] <= 3'b101;
      // memory_array[26578] <= 3'b101;
      // memory_array[26579] <= 3'b101;
      // memory_array[26580] <= 3'b101;
      // memory_array[26581] <= 3'b101;
      // memory_array[26582] <= 3'b101;
      // memory_array[26583] <= 3'b101;
      // memory_array[26584] <= 3'b101;
      // memory_array[26585] <= 3'b101;
      // memory_array[26586] <= 3'b101;
      // memory_array[26587] <= 3'b101;
      // memory_array[26588] <= 3'b101;
      // memory_array[26589] <= 3'b101;
      // memory_array[26590] <= 3'b101;
      // memory_array[26591] <= 3'b101;
      // memory_array[26592] <= 3'b111;
      // memory_array[26593] <= 3'b111;
      // memory_array[26594] <= 3'b111;
      // memory_array[26595] <= 3'b111;
      // memory_array[26596] <= 3'b111;
      // memory_array[26597] <= 3'b111;
      // memory_array[26598] <= 3'b111;
      // memory_array[26599] <= 3'b111;
      // memory_array[26600] <= 3'b111;
      // memory_array[26601] <= 3'b111;
      // memory_array[26602] <= 3'b111;
      // memory_array[26603] <= 3'b111;
      // memory_array[26604] <= 3'b111;
      // memory_array[26605] <= 3'b111;
      // memory_array[26606] <= 3'b111;
      // memory_array[26607] <= 3'b111;
      // memory_array[26608] <= 3'b101;
      // memory_array[26609] <= 3'b101;
      // memory_array[26610] <= 3'b101;
      // memory_array[26611] <= 3'b101;
      // memory_array[26612] <= 3'b101;
      // memory_array[26613] <= 3'b101;
      // memory_array[26614] <= 3'b000;
      // memory_array[26615] <= 3'b101;
      // memory_array[26616] <= 3'b000;
      // memory_array[26617] <= 3'b101;
      // memory_array[26618] <= 3'b000;
      // memory_array[26619] <= 3'b000;
      // memory_array[26620] <= 3'b101;
      // memory_array[26621] <= 3'b101;
      // memory_array[26622] <= 3'b101;
      // memory_array[26623] <= 3'b101;
      // memory_array[26624] <= 3'b101;
      // memory_array[26625] <= 3'b101;
      // memory_array[26626] <= 3'b101;
      // memory_array[26627] <= 3'b101;
      // memory_array[26628] <= 3'b101;
      // memory_array[26629] <= 3'b101;
      // memory_array[26630] <= 3'b101;
      // memory_array[26631] <= 3'b101;
      // memory_array[26632] <= 3'b101;
      // memory_array[26633] <= 3'b101;
      // memory_array[26634] <= 3'b101;
      // memory_array[26635] <= 3'b101;
      // memory_array[26636] <= 3'b101;
      // memory_array[26637] <= 3'b101;
      // memory_array[26638] <= 3'b101;
      // memory_array[26639] <= 3'b101;
      // memory_array[26640] <= 3'b101;
      // memory_array[26641] <= 3'b101;
      // memory_array[26642] <= 3'b101;
      // memory_array[26643] <= 3'b101;
      // memory_array[26644] <= 3'b101;
      // memory_array[26645] <= 3'b101;
      // memory_array[26646] <= 3'b101;
      // memory_array[26647] <= 3'b101;
      // memory_array[26648] <= 3'b101;
      // memory_array[26649] <= 3'b101;
      // memory_array[26650] <= 3'b101;
      // memory_array[26651] <= 3'b101;
      // memory_array[26652] <= 3'b101;
      // memory_array[26653] <= 3'b101;
      // memory_array[26654] <= 3'b101;
      // memory_array[26655] <= 3'b101;
      // memory_array[26656] <= 3'b101;
      // memory_array[26657] <= 3'b101;
      // memory_array[26658] <= 3'b101;
      // memory_array[26659] <= 3'b000;
      // memory_array[26660] <= 3'b101;
      // memory_array[26661] <= 3'b000;
      // memory_array[26662] <= 3'b101;
      // memory_array[26663] <= 3'b000;
      // memory_array[26664] <= 3'b000;
      // memory_array[26665] <= 3'b101;
      // memory_array[26666] <= 3'b101;
      // memory_array[26667] <= 3'b101;
      // memory_array[26668] <= 3'b101;
      // memory_array[26669] <= 3'b101;
      // memory_array[26670] <= 3'b101;
      // memory_array[26671] <= 3'b101;
      // memory_array[26672] <= 3'b101;
      // memory_array[26673] <= 3'b101;
      // memory_array[26674] <= 3'b101;
      // memory_array[26675] <= 3'b101;
      // memory_array[26676] <= 3'b101;
      // memory_array[26677] <= 3'b101;
      // memory_array[26678] <= 3'b101;
      // memory_array[26679] <= 3'b101;
      // memory_array[26680] <= 3'b101;
      // memory_array[26681] <= 3'b101;
      // memory_array[26682] <= 3'b101;
      // memory_array[26683] <= 3'b101;
      // memory_array[26684] <= 3'b101;
      // memory_array[26685] <= 3'b101;
      // memory_array[26686] <= 3'b101;
      // memory_array[26687] <= 3'b101;
      // memory_array[26688] <= 3'b101;
      // memory_array[26689] <= 3'b101;
      // memory_array[26690] <= 3'b101;
      // memory_array[26691] <= 3'b101;
      // memory_array[26692] <= 3'b101;
      // memory_array[26693] <= 3'b101;
      // memory_array[26694] <= 3'b101;
      // memory_array[26695] <= 3'b101;
      // memory_array[26696] <= 3'b101;
      // memory_array[26697] <= 3'b101;
      // memory_array[26698] <= 3'b101;
      // memory_array[26699] <= 3'b101;
      // memory_array[26700] <= 3'b101;
      // memory_array[26701] <= 3'b101;
      // memory_array[26702] <= 3'b101;
      // memory_array[26703] <= 3'b101;
      // memory_array[26704] <= 3'b101;
      // memory_array[26705] <= 3'b101;
      // memory_array[26706] <= 3'b101;
      // memory_array[26707] <= 3'b101;
      // memory_array[26708] <= 3'b101;
      // memory_array[26709] <= 3'b101;
      // memory_array[26710] <= 3'b101;
      // memory_array[26711] <= 3'b101;
      // memory_array[26712] <= 3'b101;
      // memory_array[26713] <= 3'b101;
      // memory_array[26714] <= 3'b101;
      // memory_array[26715] <= 3'b101;
      // memory_array[26716] <= 3'b101;
      // memory_array[26717] <= 3'b101;
      // memory_array[26718] <= 3'b101;
      // memory_array[26719] <= 3'b101;
      // memory_array[26720] <= 3'b101;
      // memory_array[26721] <= 3'b101;
      // memory_array[26722] <= 3'b101;
      // memory_array[26723] <= 3'b101;
      // memory_array[26724] <= 3'b101;
      // memory_array[26725] <= 3'b101;
      // memory_array[26726] <= 3'b101;
      // memory_array[26727] <= 3'b101;
      // memory_array[26728] <= 3'b101;
      // memory_array[26729] <= 3'b101;
      // memory_array[26730] <= 3'b101;
      // memory_array[26731] <= 3'b101;
      // memory_array[26732] <= 3'b101;
      // memory_array[26733] <= 3'b101;
      // memory_array[26734] <= 3'b000;
      // memory_array[26735] <= 3'b101;
      // memory_array[26736] <= 3'b000;
      // memory_array[26737] <= 3'b101;
      // memory_array[26738] <= 3'b000;
      // memory_array[26739] <= 3'b000;
      // memory_array[26740] <= 3'b101;
      // memory_array[26741] <= 3'b101;
      // memory_array[26742] <= 3'b101;
      // memory_array[26743] <= 3'b101;
      // memory_array[26744] <= 3'b101;
      // memory_array[26745] <= 3'b101;
      // memory_array[26746] <= 3'b101;
      // memory_array[26747] <= 3'b101;
      // memory_array[26748] <= 3'b101;
      // memory_array[26749] <= 3'b101;
      // memory_array[26750] <= 3'b101;
      // memory_array[26751] <= 3'b101;
      // memory_array[26752] <= 3'b101;
      // memory_array[26753] <= 3'b101;
      // memory_array[26754] <= 3'b101;
      // memory_array[26755] <= 3'b101;
      // memory_array[26756] <= 3'b101;
      // memory_array[26757] <= 3'b101;
      // memory_array[26758] <= 3'b101;
      // memory_array[26759] <= 3'b101;
      // memory_array[26760] <= 3'b101;
      // memory_array[26761] <= 3'b101;
      // memory_array[26762] <= 3'b101;
      // memory_array[26763] <= 3'b101;
      // memory_array[26764] <= 3'b101;
      // memory_array[26765] <= 3'b101;
      // memory_array[26766] <= 3'b101;
      // memory_array[26767] <= 3'b101;
      // memory_array[26768] <= 3'b101;
      // memory_array[26769] <= 3'b101;
      // memory_array[26770] <= 3'b101;
      // memory_array[26771] <= 3'b101;
      // memory_array[26772] <= 3'b101;
      // memory_array[26773] <= 3'b101;
      // memory_array[26774] <= 3'b101;
      // memory_array[26775] <= 3'b101;
      // memory_array[26776] <= 3'b101;
      // memory_array[26777] <= 3'b101;
      // memory_array[26778] <= 3'b101;
      // memory_array[26779] <= 3'b000;
      // memory_array[26780] <= 3'b101;
      // memory_array[26781] <= 3'b000;
      // memory_array[26782] <= 3'b101;
      // memory_array[26783] <= 3'b000;
      // memory_array[26784] <= 3'b000;
      // memory_array[26785] <= 3'b101;
      // memory_array[26786] <= 3'b101;
      // memory_array[26787] <= 3'b101;
      // memory_array[26788] <= 3'b101;
      // memory_array[26789] <= 3'b101;
      // memory_array[26790] <= 3'b101;
      // memory_array[26791] <= 3'b101;
      // memory_array[26792] <= 3'b111;
      // memory_array[26793] <= 3'b111;
      // memory_array[26794] <= 3'b111;
      // memory_array[26795] <= 3'b111;
      // memory_array[26796] <= 3'b111;
      // memory_array[26797] <= 3'b111;
      // memory_array[26798] <= 3'b111;
      // memory_array[26799] <= 3'b111;
      // memory_array[26800] <= 3'b111;
      // memory_array[26801] <= 3'b111;
      // memory_array[26802] <= 3'b111;
      // memory_array[26803] <= 3'b101;
      // memory_array[26804] <= 3'b101;
      // memory_array[26805] <= 3'b101;
      // memory_array[26806] <= 3'b111;
      // memory_array[26807] <= 3'b111;
      // memory_array[26808] <= 3'b101;
      // memory_array[26809] <= 3'b101;
      // memory_array[26810] <= 3'b101;
      // memory_array[26811] <= 3'b101;
      // memory_array[26812] <= 3'b000;
      // memory_array[26813] <= 3'b000;
      // memory_array[26814] <= 3'b101;
      // memory_array[26815] <= 3'b101;
      // memory_array[26816] <= 3'b101;
      // memory_array[26817] <= 3'b101;
      // memory_array[26818] <= 3'b000;
      // memory_array[26819] <= 3'b000;
      // memory_array[26820] <= 3'b101;
      // memory_array[26821] <= 3'b000;
      // memory_array[26822] <= 3'b101;
      // memory_array[26823] <= 3'b101;
      // memory_array[26824] <= 3'b101;
      // memory_array[26825] <= 3'b101;
      // memory_array[26826] <= 3'b000;
      // memory_array[26827] <= 3'b000;
      // memory_array[26828] <= 3'b000;
      // memory_array[26829] <= 3'b000;
      // memory_array[26830] <= 3'b101;
      // memory_array[26831] <= 3'b101;
      // memory_array[26832] <= 3'b111;
      // memory_array[26833] <= 3'b111;
      // memory_array[26834] <= 3'b000;
      // memory_array[26835] <= 3'b000;
      // memory_array[26836] <= 3'b000;
      // memory_array[26837] <= 3'b000;
      // memory_array[26838] <= 3'b000;
      // memory_array[26839] <= 3'b101;
      // memory_array[26840] <= 3'b000;
      // memory_array[26841] <= 3'b101;
      // memory_array[26842] <= 3'b000;
      // memory_array[26843] <= 3'b000;
      // memory_array[26844] <= 3'b000;
      // memory_array[26845] <= 3'b000;
      // memory_array[26846] <= 3'b101;
      // memory_array[26847] <= 3'b101;
      // memory_array[26848] <= 3'b000;
      // memory_array[26849] <= 3'b101;
      // memory_array[26850] <= 3'b111;
      // memory_array[26851] <= 3'b101;
      // memory_array[26852] <= 3'b101;
      // memory_array[26853] <= 3'b101;
      // memory_array[26854] <= 3'b101;
      // memory_array[26855] <= 3'b101;
      // memory_array[26856] <= 3'b101;
      // memory_array[26857] <= 3'b000;
      // memory_array[26858] <= 3'b000;
      // memory_array[26859] <= 3'b101;
      // memory_array[26860] <= 3'b101;
      // memory_array[26861] <= 3'b101;
      // memory_array[26862] <= 3'b101;
      // memory_array[26863] <= 3'b000;
      // memory_array[26864] <= 3'b000;
      // memory_array[26865] <= 3'b101;
      // memory_array[26866] <= 3'b000;
      // memory_array[26867] <= 3'b101;
      // memory_array[26868] <= 3'b101;
      // memory_array[26869] <= 3'b101;
      // memory_array[26870] <= 3'b101;
      // memory_array[26871] <= 3'b101;
      // memory_array[26872] <= 3'b101;
      // memory_array[26873] <= 3'b101;
      // memory_array[26874] <= 3'b000;
      // memory_array[26875] <= 3'b101;
      // memory_array[26876] <= 3'b101;
      // memory_array[26877] <= 3'b101;
      // memory_array[26878] <= 3'b101;
      // memory_array[26879] <= 3'b000;
      // memory_array[26880] <= 3'b000;
      // memory_array[26881] <= 3'b000;
      // memory_array[26882] <= 3'b000;
      // memory_array[26883] <= 3'b000;
      // memory_array[26884] <= 3'b101;
      // memory_array[26885] <= 3'b111;
      // memory_array[26886] <= 3'b000;
      // memory_array[26887] <= 3'b000;
      // memory_array[26888] <= 3'b000;
      // memory_array[26889] <= 3'b000;
      // memory_array[26890] <= 3'b000;
      // memory_array[26891] <= 3'b000;
      // memory_array[26892] <= 3'b101;
      // memory_array[26893] <= 3'b101;
      // memory_array[26894] <= 3'b101;
      // memory_array[26895] <= 3'b101;
      // memory_array[26896] <= 3'b000;
      // memory_array[26897] <= 3'b000;
      // memory_array[26898] <= 3'b111;
      // memory_array[26899] <= 3'b101;
      // memory_array[26900] <= 3'b101;
      // memory_array[26901] <= 3'b111;
      // memory_array[26902] <= 3'b000;
      // memory_array[26903] <= 3'b000;
      // memory_array[26904] <= 3'b000;
      // memory_array[26905] <= 3'b101;
      // memory_array[26906] <= 3'b101;
      // memory_array[26907] <= 3'b111;
      // memory_array[26908] <= 3'b111;
      // memory_array[26909] <= 3'b000;
      // memory_array[26910] <= 3'b000;
      // memory_array[26911] <= 3'b000;
      // memory_array[26912] <= 3'b000;
      // memory_array[26913] <= 3'b000;
      // memory_array[26914] <= 3'b101;
      // memory_array[26915] <= 3'b000;
      // memory_array[26916] <= 3'b101;
      // memory_array[26917] <= 3'b000;
      // memory_array[26918] <= 3'b000;
      // memory_array[26919] <= 3'b000;
      // memory_array[26920] <= 3'b000;
      // memory_array[26921] <= 3'b101;
      // memory_array[26922] <= 3'b101;
      // memory_array[26923] <= 3'b000;
      // memory_array[26924] <= 3'b101;
      // memory_array[26925] <= 3'b111;
      // memory_array[26926] <= 3'b101;
      // memory_array[26927] <= 3'b101;
      // memory_array[26928] <= 3'b101;
      // memory_array[26929] <= 3'b101;
      // memory_array[26930] <= 3'b101;
      // memory_array[26931] <= 3'b101;
      // memory_array[26932] <= 3'b000;
      // memory_array[26933] <= 3'b000;
      // memory_array[26934] <= 3'b101;
      // memory_array[26935] <= 3'b101;
      // memory_array[26936] <= 3'b101;
      // memory_array[26937] <= 3'b101;
      // memory_array[26938] <= 3'b000;
      // memory_array[26939] <= 3'b000;
      // memory_array[26940] <= 3'b101;
      // memory_array[26941] <= 3'b000;
      // memory_array[26942] <= 3'b101;
      // memory_array[26943] <= 3'b101;
      // memory_array[26944] <= 3'b101;
      // memory_array[26945] <= 3'b101;
      // memory_array[26946] <= 3'b101;
      // memory_array[26947] <= 3'b101;
      // memory_array[26948] <= 3'b101;
      // memory_array[26949] <= 3'b000;
      // memory_array[26950] <= 3'b101;
      // memory_array[26951] <= 3'b101;
      // memory_array[26952] <= 3'b101;
      // memory_array[26953] <= 3'b101;
      // memory_array[26954] <= 3'b000;
      // memory_array[26955] <= 3'b000;
      // memory_array[26956] <= 3'b000;
      // memory_array[26957] <= 3'b000;
      // memory_array[26958] <= 3'b000;
      // memory_array[26959] <= 3'b101;
      // memory_array[26960] <= 3'b111;
      // memory_array[26961] <= 3'b000;
      // memory_array[26962] <= 3'b000;
      // memory_array[26963] <= 3'b000;
      // memory_array[26964] <= 3'b000;
      // memory_array[26965] <= 3'b000;
      // memory_array[26966] <= 3'b000;
      // memory_array[26967] <= 3'b101;
      // memory_array[26968] <= 3'b101;
      // memory_array[26969] <= 3'b101;
      // memory_array[26970] <= 3'b101;
      // memory_array[26971] <= 3'b000;
      // memory_array[26972] <= 3'b000;
      // memory_array[26973] <= 3'b111;
      // memory_array[26974] <= 3'b101;
      // memory_array[26975] <= 3'b101;
      // memory_array[26976] <= 3'b101;
      // memory_array[26977] <= 3'b000;
      // memory_array[26978] <= 3'b000;
      // memory_array[26979] <= 3'b101;
      // memory_array[26980] <= 3'b101;
      // memory_array[26981] <= 3'b101;
      // memory_array[26982] <= 3'b101;
      // memory_array[26983] <= 3'b000;
      // memory_array[26984] <= 3'b000;
      // memory_array[26985] <= 3'b101;
      // memory_array[26986] <= 3'b000;
      // memory_array[26987] <= 3'b101;
      // memory_array[26988] <= 3'b101;
      // memory_array[26989] <= 3'b101;
      // memory_array[26990] <= 3'b101;
      // memory_array[26991] <= 3'b101;
      // memory_array[26992] <= 3'b111;
      // memory_array[26993] <= 3'b111;
      // memory_array[26994] <= 3'b111;
      // memory_array[26995] <= 3'b101;
      // memory_array[26996] <= 3'b101;
      // memory_array[26997] <= 3'b111;
      // memory_array[26998] <= 3'b111;
      // memory_array[26999] <= 3'b111;
      // memory_array[27000] <= 3'b111;
      // memory_array[27001] <= 3'b111;
      // memory_array[27002] <= 3'b101;
      // memory_array[27003] <= 3'b111;
      // memory_array[27004] <= 3'b101;
      // memory_array[27005] <= 3'b101;
      // memory_array[27006] <= 3'b111;
      // memory_array[27007] <= 3'b111;
      // memory_array[27008] <= 3'b101;
      // memory_array[27009] <= 3'b101;
      // memory_array[27010] <= 3'b101;
      // memory_array[27011] <= 3'b101;
      // memory_array[27012] <= 3'b101;
      // memory_array[27013] <= 3'b101;
      // memory_array[27014] <= 3'b101;
      // memory_array[27015] <= 3'b101;
      // memory_array[27016] <= 3'b000;
      // memory_array[27017] <= 3'b101;
      // memory_array[27018] <= 3'b111;
      // memory_array[27019] <= 3'b000;
      // memory_array[27020] <= 3'b000;
      // memory_array[27021] <= 3'b000;
      // memory_array[27022] <= 3'b101;
      // memory_array[27023] <= 3'b101;
      // memory_array[27024] <= 3'b101;
      // memory_array[27025] <= 3'b101;
      // memory_array[27026] <= 3'b101;
      // memory_array[27027] <= 3'b101;
      // memory_array[27028] <= 3'b101;
      // memory_array[27029] <= 3'b111;
      // memory_array[27030] <= 3'b101;
      // memory_array[27031] <= 3'b101;
      // memory_array[27032] <= 3'b000;
      // memory_array[27033] <= 3'b101;
      // memory_array[27034] <= 3'b101;
      // memory_array[27035] <= 3'b101;
      // memory_array[27036] <= 3'b101;
      // memory_array[27037] <= 3'b101;
      // memory_array[27038] <= 3'b101;
      // memory_array[27039] <= 3'b000;
      // memory_array[27040] <= 3'b101;
      // memory_array[27041] <= 3'b000;
      // memory_array[27042] <= 3'b101;
      // memory_array[27043] <= 3'b101;
      // memory_array[27044] <= 3'b101;
      // memory_array[27045] <= 3'b101;
      // memory_array[27046] <= 3'b000;
      // memory_array[27047] <= 3'b101;
      // memory_array[27048] <= 3'b101;
      // memory_array[27049] <= 3'b101;
      // memory_array[27050] <= 3'b101;
      // memory_array[27051] <= 3'b101;
      // memory_array[27052] <= 3'b101;
      // memory_array[27053] <= 3'b101;
      // memory_array[27054] <= 3'b101;
      // memory_array[27055] <= 3'b101;
      // memory_array[27056] <= 3'b101;
      // memory_array[27057] <= 3'b101;
      // memory_array[27058] <= 3'b101;
      // memory_array[27059] <= 3'b101;
      // memory_array[27060] <= 3'b101;
      // memory_array[27061] <= 3'b000;
      // memory_array[27062] <= 3'b101;
      // memory_array[27063] <= 3'b111;
      // memory_array[27064] <= 3'b000;
      // memory_array[27065] <= 3'b000;
      // memory_array[27066] <= 3'b000;
      // memory_array[27067] <= 3'b101;
      // memory_array[27068] <= 3'b101;
      // memory_array[27069] <= 3'b101;
      // memory_array[27070] <= 3'b101;
      // memory_array[27071] <= 3'b101;
      // memory_array[27072] <= 3'b101;
      // memory_array[27073] <= 3'b000;
      // memory_array[27074] <= 3'b101;
      // memory_array[27075] <= 3'b111;
      // memory_array[27076] <= 3'b111;
      // memory_array[27077] <= 3'b101;
      // memory_array[27078] <= 3'b101;
      // memory_array[27079] <= 3'b101;
      // memory_array[27080] <= 3'b101;
      // memory_array[27081] <= 3'b101;
      // memory_array[27082] <= 3'b000;
      // memory_array[27083] <= 3'b101;
      // memory_array[27084] <= 3'b101;
      // memory_array[27085] <= 3'b111;
      // memory_array[27086] <= 3'b101;
      // memory_array[27087] <= 3'b101;
      // memory_array[27088] <= 3'b101;
      // memory_array[27089] <= 3'b101;
      // memory_array[27090] <= 3'b101;
      // memory_array[27091] <= 3'b000;
      // memory_array[27092] <= 3'b000;
      // memory_array[27093] <= 3'b000;
      // memory_array[27094] <= 3'b101;
      // memory_array[27095] <= 3'b101;
      // memory_array[27096] <= 3'b101;
      // memory_array[27097] <= 3'b000;
      // memory_array[27098] <= 3'b101;
      // memory_array[27099] <= 3'b101;
      // memory_array[27100] <= 3'b101;
      // memory_array[27101] <= 3'b111;
      // memory_array[27102] <= 3'b101;
      // memory_array[27103] <= 3'b101;
      // memory_array[27104] <= 3'b111;
      // memory_array[27105] <= 3'b101;
      // memory_array[27106] <= 3'b101;
      // memory_array[27107] <= 3'b000;
      // memory_array[27108] <= 3'b101;
      // memory_array[27109] <= 3'b101;
      // memory_array[27110] <= 3'b101;
      // memory_array[27111] <= 3'b101;
      // memory_array[27112] <= 3'b101;
      // memory_array[27113] <= 3'b101;
      // memory_array[27114] <= 3'b000;
      // memory_array[27115] <= 3'b101;
      // memory_array[27116] <= 3'b000;
      // memory_array[27117] <= 3'b101;
      // memory_array[27118] <= 3'b101;
      // memory_array[27119] <= 3'b101;
      // memory_array[27120] <= 3'b101;
      // memory_array[27121] <= 3'b000;
      // memory_array[27122] <= 3'b101;
      // memory_array[27123] <= 3'b101;
      // memory_array[27124] <= 3'b101;
      // memory_array[27125] <= 3'b101;
      // memory_array[27126] <= 3'b101;
      // memory_array[27127] <= 3'b101;
      // memory_array[27128] <= 3'b101;
      // memory_array[27129] <= 3'b101;
      // memory_array[27130] <= 3'b101;
      // memory_array[27131] <= 3'b101;
      // memory_array[27132] <= 3'b101;
      // memory_array[27133] <= 3'b101;
      // memory_array[27134] <= 3'b101;
      // memory_array[27135] <= 3'b101;
      // memory_array[27136] <= 3'b000;
      // memory_array[27137] <= 3'b101;
      // memory_array[27138] <= 3'b111;
      // memory_array[27139] <= 3'b000;
      // memory_array[27140] <= 3'b000;
      // memory_array[27141] <= 3'b000;
      // memory_array[27142] <= 3'b101;
      // memory_array[27143] <= 3'b101;
      // memory_array[27144] <= 3'b101;
      // memory_array[27145] <= 3'b101;
      // memory_array[27146] <= 3'b101;
      // memory_array[27147] <= 3'b101;
      // memory_array[27148] <= 3'b000;
      // memory_array[27149] <= 3'b101;
      // memory_array[27150] <= 3'b111;
      // memory_array[27151] <= 3'b111;
      // memory_array[27152] <= 3'b101;
      // memory_array[27153] <= 3'b101;
      // memory_array[27154] <= 3'b101;
      // memory_array[27155] <= 3'b101;
      // memory_array[27156] <= 3'b101;
      // memory_array[27157] <= 3'b000;
      // memory_array[27158] <= 3'b101;
      // memory_array[27159] <= 3'b101;
      // memory_array[27160] <= 3'b111;
      // memory_array[27161] <= 3'b101;
      // memory_array[27162] <= 3'b101;
      // memory_array[27163] <= 3'b101;
      // memory_array[27164] <= 3'b101;
      // memory_array[27165] <= 3'b101;
      // memory_array[27166] <= 3'b000;
      // memory_array[27167] <= 3'b000;
      // memory_array[27168] <= 3'b000;
      // memory_array[27169] <= 3'b101;
      // memory_array[27170] <= 3'b101;
      // memory_array[27171] <= 3'b101;
      // memory_array[27172] <= 3'b000;
      // memory_array[27173] <= 3'b101;
      // memory_array[27174] <= 3'b101;
      // memory_array[27175] <= 3'b101;
      // memory_array[27176] <= 3'b101;
      // memory_array[27177] <= 3'b101;
      // memory_array[27178] <= 3'b101;
      // memory_array[27179] <= 3'b101;
      // memory_array[27180] <= 3'b101;
      // memory_array[27181] <= 3'b000;
      // memory_array[27182] <= 3'b101;
      // memory_array[27183] <= 3'b111;
      // memory_array[27184] <= 3'b000;
      // memory_array[27185] <= 3'b000;
      // memory_array[27186] <= 3'b000;
      // memory_array[27187] <= 3'b101;
      // memory_array[27188] <= 3'b101;
      // memory_array[27189] <= 3'b101;
      // memory_array[27190] <= 3'b101;
      // memory_array[27191] <= 3'b101;
      // memory_array[27192] <= 3'b111;
      // memory_array[27193] <= 3'b111;
      // memory_array[27194] <= 3'b111;
      // memory_array[27195] <= 3'b101;
      // memory_array[27196] <= 3'b101;
      // memory_array[27197] <= 3'b111;
      // memory_array[27198] <= 3'b111;
      // memory_array[27199] <= 3'b111;
      // memory_array[27200] <= 3'b111;
      // memory_array[27201] <= 3'b111;
      // memory_array[27202] <= 3'b111;
      // memory_array[27203] <= 3'b111;
      // memory_array[27204] <= 3'b111;
      // memory_array[27205] <= 3'b101;
      // memory_array[27206] <= 3'b101;
      // memory_array[27207] <= 3'b111;
      // memory_array[27208] <= 3'b101;
      // memory_array[27209] <= 3'b101;
      // memory_array[27210] <= 3'b101;
      // memory_array[27211] <= 3'b101;
      // memory_array[27212] <= 3'b000;
      // memory_array[27213] <= 3'b101;
      // memory_array[27214] <= 3'b101;
      // memory_array[27215] <= 3'b111;
      // memory_array[27216] <= 3'b000;
      // memory_array[27217] <= 3'b000;
      // memory_array[27218] <= 3'b101;
      // memory_array[27219] <= 3'b000;
      // memory_array[27220] <= 3'b101;
      // memory_array[27221] <= 3'b101;
      // memory_array[27222] <= 3'b101;
      // memory_array[27223] <= 3'b101;
      // memory_array[27224] <= 3'b101;
      // memory_array[27225] <= 3'b101;
      // memory_array[27226] <= 3'b101;
      // memory_array[27227] <= 3'b101;
      // memory_array[27228] <= 3'b101;
      // memory_array[27229] <= 3'b111;
      // memory_array[27230] <= 3'b111;
      // memory_array[27231] <= 3'b101;
      // memory_array[27232] <= 3'b101;
      // memory_array[27233] <= 3'b101;
      // memory_array[27234] <= 3'b101;
      // memory_array[27235] <= 3'b101;
      // memory_array[27236] <= 3'b101;
      // memory_array[27237] <= 3'b101;
      // memory_array[27238] <= 3'b101;
      // memory_array[27239] <= 3'b000;
      // memory_array[27240] <= 3'b000;
      // memory_array[27241] <= 3'b101;
      // memory_array[27242] <= 3'b101;
      // memory_array[27243] <= 3'b111;
      // memory_array[27244] <= 3'b101;
      // memory_array[27245] <= 3'b101;
      // memory_array[27246] <= 3'b000;
      // memory_array[27247] <= 3'b000;
      // memory_array[27248] <= 3'b000;
      // memory_array[27249] <= 3'b101;
      // memory_array[27250] <= 3'b101;
      // memory_array[27251] <= 3'b101;
      // memory_array[27252] <= 3'b101;
      // memory_array[27253] <= 3'b101;
      // memory_array[27254] <= 3'b101;
      // memory_array[27255] <= 3'b101;
      // memory_array[27256] <= 3'b101;
      // memory_array[27257] <= 3'b000;
      // memory_array[27258] <= 3'b101;
      // memory_array[27259] <= 3'b101;
      // memory_array[27260] <= 3'b111;
      // memory_array[27261] <= 3'b000;
      // memory_array[27262] <= 3'b000;
      // memory_array[27263] <= 3'b101;
      // memory_array[27264] <= 3'b000;
      // memory_array[27265] <= 3'b101;
      // memory_array[27266] <= 3'b101;
      // memory_array[27267] <= 3'b101;
      // memory_array[27268] <= 3'b101;
      // memory_array[27269] <= 3'b101;
      // memory_array[27270] <= 3'b101;
      // memory_array[27271] <= 3'b101;
      // memory_array[27272] <= 3'b000;
      // memory_array[27273] <= 3'b000;
      // memory_array[27274] <= 3'b101;
      // memory_array[27275] <= 3'b101;
      // memory_array[27276] <= 3'b000;
      // memory_array[27277] <= 3'b000;
      // memory_array[27278] <= 3'b101;
      // memory_array[27279] <= 3'b101;
      // memory_array[27280] <= 3'b101;
      // memory_array[27281] <= 3'b000;
      // memory_array[27282] <= 3'b111;
      // memory_array[27283] <= 3'b101;
      // memory_array[27284] <= 3'b101;
      // memory_array[27285] <= 3'b101;
      // memory_array[27286] <= 3'b101;
      // memory_array[27287] <= 3'b101;
      // memory_array[27288] <= 3'b101;
      // memory_array[27289] <= 3'b101;
      // memory_array[27290] <= 3'b101;
      // memory_array[27291] <= 3'b101;
      // memory_array[27292] <= 3'b101;
      // memory_array[27293] <= 3'b000;
      // memory_array[27294] <= 3'b111;
      // memory_array[27295] <= 3'b111;
      // memory_array[27296] <= 3'b101;
      // memory_array[27297] <= 3'b000;
      // memory_array[27298] <= 3'b101;
      // memory_array[27299] <= 3'b101;
      // memory_array[27300] <= 3'b101;
      // memory_array[27301] <= 3'b111;
      // memory_array[27302] <= 3'b101;
      // memory_array[27303] <= 3'b101;
      // memory_array[27304] <= 3'b111;
      // memory_array[27305] <= 3'b111;
      // memory_array[27306] <= 3'b101;
      // memory_array[27307] <= 3'b101;
      // memory_array[27308] <= 3'b101;
      // memory_array[27309] <= 3'b101;
      // memory_array[27310] <= 3'b101;
      // memory_array[27311] <= 3'b101;
      // memory_array[27312] <= 3'b101;
      // memory_array[27313] <= 3'b101;
      // memory_array[27314] <= 3'b000;
      // memory_array[27315] <= 3'b000;
      // memory_array[27316] <= 3'b101;
      // memory_array[27317] <= 3'b101;
      // memory_array[27318] <= 3'b111;
      // memory_array[27319] <= 3'b101;
      // memory_array[27320] <= 3'b101;
      // memory_array[27321] <= 3'b000;
      // memory_array[27322] <= 3'b000;
      // memory_array[27323] <= 3'b000;
      // memory_array[27324] <= 3'b101;
      // memory_array[27325] <= 3'b101;
      // memory_array[27326] <= 3'b101;
      // memory_array[27327] <= 3'b101;
      // memory_array[27328] <= 3'b101;
      // memory_array[27329] <= 3'b101;
      // memory_array[27330] <= 3'b101;
      // memory_array[27331] <= 3'b101;
      // memory_array[27332] <= 3'b000;
      // memory_array[27333] <= 3'b101;
      // memory_array[27334] <= 3'b101;
      // memory_array[27335] <= 3'b111;
      // memory_array[27336] <= 3'b000;
      // memory_array[27337] <= 3'b000;
      // memory_array[27338] <= 3'b101;
      // memory_array[27339] <= 3'b000;
      // memory_array[27340] <= 3'b101;
      // memory_array[27341] <= 3'b101;
      // memory_array[27342] <= 3'b101;
      // memory_array[27343] <= 3'b101;
      // memory_array[27344] <= 3'b101;
      // memory_array[27345] <= 3'b101;
      // memory_array[27346] <= 3'b101;
      // memory_array[27347] <= 3'b000;
      // memory_array[27348] <= 3'b000;
      // memory_array[27349] <= 3'b101;
      // memory_array[27350] <= 3'b101;
      // memory_array[27351] <= 3'b000;
      // memory_array[27352] <= 3'b000;
      // memory_array[27353] <= 3'b101;
      // memory_array[27354] <= 3'b101;
      // memory_array[27355] <= 3'b101;
      // memory_array[27356] <= 3'b000;
      // memory_array[27357] <= 3'b111;
      // memory_array[27358] <= 3'b101;
      // memory_array[27359] <= 3'b101;
      // memory_array[27360] <= 3'b101;
      // memory_array[27361] <= 3'b101;
      // memory_array[27362] <= 3'b101;
      // memory_array[27363] <= 3'b101;
      // memory_array[27364] <= 3'b101;
      // memory_array[27365] <= 3'b101;
      // memory_array[27366] <= 3'b101;
      // memory_array[27367] <= 3'b101;
      // memory_array[27368] <= 3'b000;
      // memory_array[27369] <= 3'b111;
      // memory_array[27370] <= 3'b111;
      // memory_array[27371] <= 3'b101;
      // memory_array[27372] <= 3'b000;
      // memory_array[27373] <= 3'b101;
      // memory_array[27374] <= 3'b101;
      // memory_array[27375] <= 3'b101;
      // memory_array[27376] <= 3'b101;
      // memory_array[27377] <= 3'b000;
      // memory_array[27378] <= 3'b101;
      // memory_array[27379] <= 3'b101;
      // memory_array[27380] <= 3'b111;
      // memory_array[27381] <= 3'b000;
      // memory_array[27382] <= 3'b000;
      // memory_array[27383] <= 3'b101;
      // memory_array[27384] <= 3'b000;
      // memory_array[27385] <= 3'b101;
      // memory_array[27386] <= 3'b101;
      // memory_array[27387] <= 3'b101;
      // memory_array[27388] <= 3'b101;
      // memory_array[27389] <= 3'b101;
      // memory_array[27390] <= 3'b101;
      // memory_array[27391] <= 3'b101;
      // memory_array[27392] <= 3'b111;
      // memory_array[27393] <= 3'b101;
      // memory_array[27394] <= 3'b101;
      // memory_array[27395] <= 3'b111;
      // memory_array[27396] <= 3'b111;
      // memory_array[27397] <= 3'b101;
      // memory_array[27398] <= 3'b101;
      // memory_array[27399] <= 3'b111;
      // memory_array[27400] <= 3'b111;
      // memory_array[27401] <= 3'b101;
      // memory_array[27402] <= 3'b101;
      // memory_array[27403] <= 3'b111;
      // memory_array[27404] <= 3'b111;
      // memory_array[27405] <= 3'b111;
      // memory_array[27406] <= 3'b101;
      // memory_array[27407] <= 3'b111;
      // memory_array[27408] <= 3'b101;
      // memory_array[27409] <= 3'b101;
      // memory_array[27410] <= 3'b101;
      // memory_array[27411] <= 3'b000;
      // memory_array[27412] <= 3'b000;
      // memory_array[27413] <= 3'b101;
      // memory_array[27414] <= 3'b111;
      // memory_array[27415] <= 3'b000;
      // memory_array[27416] <= 3'b101;
      // memory_array[27417] <= 3'b000;
      // memory_array[27418] <= 3'b111;
      // memory_array[27419] <= 3'b000;
      // memory_array[27420] <= 3'b000;
      // memory_array[27421] <= 3'b101;
      // memory_array[27422] <= 3'b000;
      // memory_array[27423] <= 3'b000;
      // memory_array[27424] <= 3'b101;
      // memory_array[27425] <= 3'b101;
      // memory_array[27426] <= 3'b101;
      // memory_array[27427] <= 3'b101;
      // memory_array[27428] <= 3'b101;
      // memory_array[27429] <= 3'b000;
      // memory_array[27430] <= 3'b000;
      // memory_array[27431] <= 3'b101;
      // memory_array[27432] <= 3'b101;
      // memory_array[27433] <= 3'b101;
      // memory_array[27434] <= 3'b101;
      // memory_array[27435] <= 3'b101;
      // memory_array[27436] <= 3'b101;
      // memory_array[27437] <= 3'b101;
      // memory_array[27438] <= 3'b101;
      // memory_array[27439] <= 3'b101;
      // memory_array[27440] <= 3'b000;
      // memory_array[27441] <= 3'b111;
      // memory_array[27442] <= 3'b101;
      // memory_array[27443] <= 3'b101;
      // memory_array[27444] <= 3'b101;
      // memory_array[27445] <= 3'b101;
      // memory_array[27446] <= 3'b101;
      // memory_array[27447] <= 3'b111;
      // memory_array[27448] <= 3'b111;
      // memory_array[27449] <= 3'b101;
      // memory_array[27450] <= 3'b101;
      // memory_array[27451] <= 3'b000;
      // memory_array[27452] <= 3'b111;
      // memory_array[27453] <= 3'b111;
      // memory_array[27454] <= 3'b101;
      // memory_array[27455] <= 3'b101;
      // memory_array[27456] <= 3'b000;
      // memory_array[27457] <= 3'b000;
      // memory_array[27458] <= 3'b101;
      // memory_array[27459] <= 3'b111;
      // memory_array[27460] <= 3'b000;
      // memory_array[27461] <= 3'b101;
      // memory_array[27462] <= 3'b000;
      // memory_array[27463] <= 3'b111;
      // memory_array[27464] <= 3'b000;
      // memory_array[27465] <= 3'b000;
      // memory_array[27466] <= 3'b101;
      // memory_array[27467] <= 3'b000;
      // memory_array[27468] <= 3'b000;
      // memory_array[27469] <= 3'b101;
      // memory_array[27470] <= 3'b101;
      // memory_array[27471] <= 3'b000;
      // memory_array[27472] <= 3'b101;
      // memory_array[27473] <= 3'b000;
      // memory_array[27474] <= 3'b101;
      // memory_array[27475] <= 3'b101;
      // memory_array[27476] <= 3'b101;
      // memory_array[27477] <= 3'b111;
      // memory_array[27478] <= 3'b111;
      // memory_array[27479] <= 3'b101;
      // memory_array[27480] <= 3'b101;
      // memory_array[27481] <= 3'b101;
      // memory_array[27482] <= 3'b000;
      // memory_array[27483] <= 3'b111;
      // memory_array[27484] <= 3'b101;
      // memory_array[27485] <= 3'b101;
      // memory_array[27486] <= 3'b000;
      // memory_array[27487] <= 3'b101;
      // memory_array[27488] <= 3'b111;
      // memory_array[27489] <= 3'b111;
      // memory_array[27490] <= 3'b111;
      // memory_array[27491] <= 3'b101;
      // memory_array[27492] <= 3'b101;
      // memory_array[27493] <= 3'b101;
      // memory_array[27494] <= 3'b000;
      // memory_array[27495] <= 3'b101;
      // memory_array[27496] <= 3'b101;
      // memory_array[27497] <= 3'b111;
      // memory_array[27498] <= 3'b101;
      // memory_array[27499] <= 3'b101;
      // memory_array[27500] <= 3'b101;
      // memory_array[27501] <= 3'b111;
      // memory_array[27502] <= 3'b101;
      // memory_array[27503] <= 3'b101;
      // memory_array[27504] <= 3'b000;
      // memory_array[27505] <= 3'b000;
      // memory_array[27506] <= 3'b101;
      // memory_array[27507] <= 3'b101;
      // memory_array[27508] <= 3'b101;
      // memory_array[27509] <= 3'b101;
      // memory_array[27510] <= 3'b101;
      // memory_array[27511] <= 3'b101;
      // memory_array[27512] <= 3'b101;
      // memory_array[27513] <= 3'b101;
      // memory_array[27514] <= 3'b101;
      // memory_array[27515] <= 3'b000;
      // memory_array[27516] <= 3'b111;
      // memory_array[27517] <= 3'b101;
      // memory_array[27518] <= 3'b101;
      // memory_array[27519] <= 3'b101;
      // memory_array[27520] <= 3'b101;
      // memory_array[27521] <= 3'b101;
      // memory_array[27522] <= 3'b111;
      // memory_array[27523] <= 3'b111;
      // memory_array[27524] <= 3'b101;
      // memory_array[27525] <= 3'b101;
      // memory_array[27526] <= 3'b000;
      // memory_array[27527] <= 3'b111;
      // memory_array[27528] <= 3'b111;
      // memory_array[27529] <= 3'b101;
      // memory_array[27530] <= 3'b101;
      // memory_array[27531] <= 3'b000;
      // memory_array[27532] <= 3'b000;
      // memory_array[27533] <= 3'b101;
      // memory_array[27534] <= 3'b111;
      // memory_array[27535] <= 3'b000;
      // memory_array[27536] <= 3'b101;
      // memory_array[27537] <= 3'b000;
      // memory_array[27538] <= 3'b111;
      // memory_array[27539] <= 3'b000;
      // memory_array[27540] <= 3'b000;
      // memory_array[27541] <= 3'b101;
      // memory_array[27542] <= 3'b000;
      // memory_array[27543] <= 3'b000;
      // memory_array[27544] <= 3'b101;
      // memory_array[27545] <= 3'b101;
      // memory_array[27546] <= 3'b000;
      // memory_array[27547] <= 3'b101;
      // memory_array[27548] <= 3'b000;
      // memory_array[27549] <= 3'b101;
      // memory_array[27550] <= 3'b101;
      // memory_array[27551] <= 3'b101;
      // memory_array[27552] <= 3'b111;
      // memory_array[27553] <= 3'b111;
      // memory_array[27554] <= 3'b101;
      // memory_array[27555] <= 3'b101;
      // memory_array[27556] <= 3'b101;
      // memory_array[27557] <= 3'b000;
      // memory_array[27558] <= 3'b111;
      // memory_array[27559] <= 3'b101;
      // memory_array[27560] <= 3'b101;
      // memory_array[27561] <= 3'b000;
      // memory_array[27562] <= 3'b101;
      // memory_array[27563] <= 3'b111;
      // memory_array[27564] <= 3'b111;
      // memory_array[27565] <= 3'b111;
      // memory_array[27566] <= 3'b101;
      // memory_array[27567] <= 3'b101;
      // memory_array[27568] <= 3'b101;
      // memory_array[27569] <= 3'b000;
      // memory_array[27570] <= 3'b101;
      // memory_array[27571] <= 3'b101;
      // memory_array[27572] <= 3'b111;
      // memory_array[27573] <= 3'b101;
      // memory_array[27574] <= 3'b101;
      // memory_array[27575] <= 3'b101;
      // memory_array[27576] <= 3'b111;
      // memory_array[27577] <= 3'b000;
      // memory_array[27578] <= 3'b101;
      // memory_array[27579] <= 3'b111;
      // memory_array[27580] <= 3'b000;
      // memory_array[27581] <= 3'b101;
      // memory_array[27582] <= 3'b000;
      // memory_array[27583] <= 3'b111;
      // memory_array[27584] <= 3'b000;
      // memory_array[27585] <= 3'b000;
      // memory_array[27586] <= 3'b101;
      // memory_array[27587] <= 3'b000;
      // memory_array[27588] <= 3'b000;
      // memory_array[27589] <= 3'b101;
      // memory_array[27590] <= 3'b101;
      // memory_array[27591] <= 3'b101;
      // memory_array[27592] <= 3'b111;
      // memory_array[27593] <= 3'b101;
      // memory_array[27594] <= 3'b101;
      // memory_array[27595] <= 3'b111;
      // memory_array[27596] <= 3'b111;
      // memory_array[27597] <= 3'b101;
      // memory_array[27598] <= 3'b101;
      // memory_array[27599] <= 3'b111;
      // memory_array[27600] <= 3'b111;
      // memory_array[27601] <= 3'b111;
      // memory_array[27602] <= 3'b111;
      // memory_array[27603] <= 3'b111;
      // memory_array[27604] <= 3'b111;
      // memory_array[27605] <= 3'b111;
      // memory_array[27606] <= 3'b111;
      // memory_array[27607] <= 3'b111;
      // memory_array[27608] <= 3'b101;
      // memory_array[27609] <= 3'b101;
      // memory_array[27610] <= 3'b000;
      // memory_array[27611] <= 3'b101;
      // memory_array[27612] <= 3'b000;
      // memory_array[27613] <= 3'b101;
      // memory_array[27614] <= 3'b101;
      // memory_array[27615] <= 3'b101;
      // memory_array[27616] <= 3'b000;
      // memory_array[27617] <= 3'b101;
      // memory_array[27618] <= 3'b000;
      // memory_array[27619] <= 3'b101;
      // memory_array[27620] <= 3'b101;
      // memory_array[27621] <= 3'b000;
      // memory_array[27622] <= 3'b101;
      // memory_array[27623] <= 3'b000;
      // memory_array[27624] <= 3'b111;
      // memory_array[27625] <= 3'b101;
      // memory_array[27626] <= 3'b101;
      // memory_array[27627] <= 3'b101;
      // memory_array[27628] <= 3'b101;
      // memory_array[27629] <= 3'b101;
      // memory_array[27630] <= 3'b101;
      // memory_array[27631] <= 3'b000;
      // memory_array[27632] <= 3'b000;
      // memory_array[27633] <= 3'b000;
      // memory_array[27634] <= 3'b000;
      // memory_array[27635] <= 3'b000;
      // memory_array[27636] <= 3'b000;
      // memory_array[27637] <= 3'b000;
      // memory_array[27638] <= 3'b101;
      // memory_array[27639] <= 3'b000;
      // memory_array[27640] <= 3'b000;
      // memory_array[27641] <= 3'b000;
      // memory_array[27642] <= 3'b101;
      // memory_array[27643] <= 3'b000;
      // memory_array[27644] <= 3'b101;
      // memory_array[27645] <= 3'b101;
      // memory_array[27646] <= 3'b000;
      // memory_array[27647] <= 3'b000;
      // memory_array[27648] <= 3'b111;
      // memory_array[27649] <= 3'b000;
      // memory_array[27650] <= 3'b000;
      // memory_array[27651] <= 3'b101;
      // memory_array[27652] <= 3'b000;
      // memory_array[27653] <= 3'b101;
      // memory_array[27654] <= 3'b101;
      // memory_array[27655] <= 3'b000;
      // memory_array[27656] <= 3'b101;
      // memory_array[27657] <= 3'b000;
      // memory_array[27658] <= 3'b101;
      // memory_array[27659] <= 3'b101;
      // memory_array[27660] <= 3'b101;
      // memory_array[27661] <= 3'b000;
      // memory_array[27662] <= 3'b000;
      // memory_array[27663] <= 3'b111;
      // memory_array[27664] <= 3'b000;
      // memory_array[27665] <= 3'b101;
      // memory_array[27666] <= 3'b000;
      // memory_array[27667] <= 3'b101;
      // memory_array[27668] <= 3'b000;
      // memory_array[27669] <= 3'b000;
      // memory_array[27670] <= 3'b000;
      // memory_array[27671] <= 3'b000;
      // memory_array[27672] <= 3'b101;
      // memory_array[27673] <= 3'b101;
      // memory_array[27674] <= 3'b000;
      // memory_array[27675] <= 3'b000;
      // memory_array[27676] <= 3'b000;
      // memory_array[27677] <= 3'b000;
      // memory_array[27678] <= 3'b000;
      // memory_array[27679] <= 3'b000;
      // memory_array[27680] <= 3'b000;
      // memory_array[27681] <= 3'b101;
      // memory_array[27682] <= 3'b000;
      // memory_array[27683] <= 3'b000;
      // memory_array[27684] <= 3'b101;
      // memory_array[27685] <= 3'b101;
      // memory_array[27686] <= 3'b000;
      // memory_array[27687] <= 3'b000;
      // memory_array[27688] <= 3'b000;
      // memory_array[27689] <= 3'b000;
      // memory_array[27690] <= 3'b000;
      // memory_array[27691] <= 3'b000;
      // memory_array[27692] <= 3'b000;
      // memory_array[27693] <= 3'b000;
      // memory_array[27694] <= 3'b000;
      // memory_array[27695] <= 3'b000;
      // memory_array[27696] <= 3'b000;
      // memory_array[27697] <= 3'b111;
      // memory_array[27698] <= 3'b101;
      // memory_array[27699] <= 3'b101;
      // memory_array[27700] <= 3'b101;
      // memory_array[27701] <= 3'b000;
      // memory_array[27702] <= 3'b000;
      // memory_array[27703] <= 3'b000;
      // memory_array[27704] <= 3'b101;
      // memory_array[27705] <= 3'b101;
      // memory_array[27706] <= 3'b000;
      // memory_array[27707] <= 3'b000;
      // memory_array[27708] <= 3'b000;
      // memory_array[27709] <= 3'b000;
      // memory_array[27710] <= 3'b000;
      // memory_array[27711] <= 3'b000;
      // memory_array[27712] <= 3'b000;
      // memory_array[27713] <= 3'b101;
      // memory_array[27714] <= 3'b000;
      // memory_array[27715] <= 3'b101;
      // memory_array[27716] <= 3'b000;
      // memory_array[27717] <= 3'b000;
      // memory_array[27718] <= 3'b000;
      // memory_array[27719] <= 3'b101;
      // memory_array[27720] <= 3'b101;
      // memory_array[27721] <= 3'b000;
      // memory_array[27722] <= 3'b000;
      // memory_array[27723] <= 3'b111;
      // memory_array[27724] <= 3'b000;
      // memory_array[27725] <= 3'b000;
      // memory_array[27726] <= 3'b101;
      // memory_array[27727] <= 3'b000;
      // memory_array[27728] <= 3'b101;
      // memory_array[27729] <= 3'b101;
      // memory_array[27730] <= 3'b000;
      // memory_array[27731] <= 3'b101;
      // memory_array[27732] <= 3'b000;
      // memory_array[27733] <= 3'b000;
      // memory_array[27734] <= 3'b000;
      // memory_array[27735] <= 3'b101;
      // memory_array[27736] <= 3'b000;
      // memory_array[27737] <= 3'b101;
      // memory_array[27738] <= 3'b000;
      // memory_array[27739] <= 3'b000;
      // memory_array[27740] <= 3'b000;
      // memory_array[27741] <= 3'b000;
      // memory_array[27742] <= 3'b101;
      // memory_array[27743] <= 3'b000;
      // memory_array[27744] <= 3'b111;
      // memory_array[27745] <= 3'b101;
      // memory_array[27746] <= 3'b000;
      // memory_array[27747] <= 3'b101;
      // memory_array[27748] <= 3'b101;
      // memory_array[27749] <= 3'b000;
      // memory_array[27750] <= 3'b000;
      // memory_array[27751] <= 3'b000;
      // memory_array[27752] <= 3'b000;
      // memory_array[27753] <= 3'b000;
      // memory_array[27754] <= 3'b000;
      // memory_array[27755] <= 3'b000;
      // memory_array[27756] <= 3'b101;
      // memory_array[27757] <= 3'b000;
      // memory_array[27758] <= 3'b000;
      // memory_array[27759] <= 3'b101;
      // memory_array[27760] <= 3'b101;
      // memory_array[27761] <= 3'b101;
      // memory_array[27762] <= 3'b000;
      // memory_array[27763] <= 3'b000;
      // memory_array[27764] <= 3'b000;
      // memory_array[27765] <= 3'b000;
      // memory_array[27766] <= 3'b000;
      // memory_array[27767] <= 3'b000;
      // memory_array[27768] <= 3'b000;
      // memory_array[27769] <= 3'b101;
      // memory_array[27770] <= 3'b101;
      // memory_array[27771] <= 3'b111;
      // memory_array[27772] <= 3'b111;
      // memory_array[27773] <= 3'b101;
      // memory_array[27774] <= 3'b101;
      // memory_array[27775] <= 3'b000;
      // memory_array[27776] <= 3'b101;
      // memory_array[27777] <= 3'b000;
      // memory_array[27778] <= 3'b101;
      // memory_array[27779] <= 3'b101;
      // memory_array[27780] <= 3'b101;
      // memory_array[27781] <= 3'b000;
      // memory_array[27782] <= 3'b101;
      // memory_array[27783] <= 3'b000;
      // memory_array[27784] <= 3'b101;
      // memory_array[27785] <= 3'b101;
      // memory_array[27786] <= 3'b000;
      // memory_array[27787] <= 3'b101;
      // memory_array[27788] <= 3'b000;
      // memory_array[27789] <= 3'b111;
      // memory_array[27790] <= 3'b101;
      // memory_array[27791] <= 3'b101;
      // memory_array[27792] <= 3'b111;
      // memory_array[27793] <= 3'b111;
      // memory_array[27794] <= 3'b111;
      // memory_array[27795] <= 3'b101;
      // memory_array[27796] <= 3'b101;
      // memory_array[27797] <= 3'b111;
      // memory_array[27798] <= 3'b111;
      // memory_array[27799] <= 3'b111;
      // memory_array[27800] <= 3'b111;
      // memory_array[27801] <= 3'b111;
      // memory_array[27802] <= 3'b101;
      // memory_array[27803] <= 3'b101;
      // memory_array[27804] <= 3'b111;
      // memory_array[27805] <= 3'b111;
      // memory_array[27806] <= 3'b111;
      // memory_array[27807] <= 3'b111;
      // memory_array[27808] <= 3'b101;
      // memory_array[27809] <= 3'b101;
      // memory_array[27810] <= 3'b000;
      // memory_array[27811] <= 3'b101;
      // memory_array[27812] <= 3'b000;
      // memory_array[27813] <= 3'b101;
      // memory_array[27814] <= 3'b111;
      // memory_array[27815] <= 3'b111;
      // memory_array[27816] <= 3'b101;
      // memory_array[27817] <= 3'b101;
      // memory_array[27818] <= 3'b000;
      // memory_array[27819] <= 3'b101;
      // memory_array[27820] <= 3'b101;
      // memory_array[27821] <= 3'b000;
      // memory_array[27822] <= 3'b000;
      // memory_array[27823] <= 3'b111;
      // memory_array[27824] <= 3'b101;
      // memory_array[27825] <= 3'b101;
      // memory_array[27826] <= 3'b101;
      // memory_array[27827] <= 3'b000;
      // memory_array[27828] <= 3'b000;
      // memory_array[27829] <= 3'b000;
      // memory_array[27830] <= 3'b101;
      // memory_array[27831] <= 3'b111;
      // memory_array[27832] <= 3'b000;
      // memory_array[27833] <= 3'b000;
      // memory_array[27834] <= 3'b111;
      // memory_array[27835] <= 3'b111;
      // memory_array[27836] <= 3'b101;
      // memory_array[27837] <= 3'b000;
      // memory_array[27838] <= 3'b111;
      // memory_array[27839] <= 3'b000;
      // memory_array[27840] <= 3'b000;
      // memory_array[27841] <= 3'b000;
      // memory_array[27842] <= 3'b000;
      // memory_array[27843] <= 3'b000;
      // memory_array[27844] <= 3'b000;
      // memory_array[27845] <= 3'b101;
      // memory_array[27846] <= 3'b000;
      // memory_array[27847] <= 3'b000;
      // memory_array[27848] <= 3'b000;
      // memory_array[27849] <= 3'b000;
      // memory_array[27850] <= 3'b101;
      // memory_array[27851] <= 3'b000;
      // memory_array[27852] <= 3'b000;
      // memory_array[27853] <= 3'b000;
      // memory_array[27854] <= 3'b000;
      // memory_array[27855] <= 3'b000;
      // memory_array[27856] <= 3'b000;
      // memory_array[27857] <= 3'b000;
      // memory_array[27858] <= 3'b000;
      // memory_array[27859] <= 3'b111;
      // memory_array[27860] <= 3'b000;
      // memory_array[27861] <= 3'b000;
      // memory_array[27862] <= 3'b000;
      // memory_array[27863] <= 3'b000;
      // memory_array[27864] <= 3'b000;
      // memory_array[27865] <= 3'b101;
      // memory_array[27866] <= 3'b000;
      // memory_array[27867] <= 3'b000;
      // memory_array[27868] <= 3'b111;
      // memory_array[27869] <= 3'b000;
      // memory_array[27870] <= 3'b000;
      // memory_array[27871] <= 3'b111;
      // memory_array[27872] <= 3'b000;
      // memory_array[27873] <= 3'b000;
      // memory_array[27874] <= 3'b000;
      // memory_array[27875] <= 3'b000;
      // memory_array[27876] <= 3'b111;
      // memory_array[27877] <= 3'b000;
      // memory_array[27878] <= 3'b000;
      // memory_array[27879] <= 3'b101;
      // memory_array[27880] <= 3'b111;
      // memory_array[27881] <= 3'b000;
      // memory_array[27882] <= 3'b111;
      // memory_array[27883] <= 3'b111;
      // memory_array[27884] <= 3'b000;
      // memory_array[27885] <= 3'b111;
      // memory_array[27886] <= 3'b000;
      // memory_array[27887] <= 3'b111;
      // memory_array[27888] <= 3'b111;
      // memory_array[27889] <= 3'b111;
      // memory_array[27890] <= 3'b111;
      // memory_array[27891] <= 3'b000;
      // memory_array[27892] <= 3'b111;
      // memory_array[27893] <= 3'b000;
      // memory_array[27894] <= 3'b111;
      // memory_array[27895] <= 3'b000;
      // memory_array[27896] <= 3'b111;
      // memory_array[27897] <= 3'b000;
      // memory_array[27898] <= 3'b101;
      // memory_array[27899] <= 3'b101;
      // memory_array[27900] <= 3'b101;
      // memory_array[27901] <= 3'b000;
      // memory_array[27902] <= 3'b111;
      // memory_array[27903] <= 3'b000;
      // memory_array[27904] <= 3'b000;
      // memory_array[27905] <= 3'b000;
      // memory_array[27906] <= 3'b000;
      // memory_array[27907] <= 3'b101;
      // memory_array[27908] <= 3'b000;
      // memory_array[27909] <= 3'b000;
      // memory_array[27910] <= 3'b000;
      // memory_array[27911] <= 3'b000;
      // memory_array[27912] <= 3'b000;
      // memory_array[27913] <= 3'b000;
      // memory_array[27914] <= 3'b101;
      // memory_array[27915] <= 3'b000;
      // memory_array[27916] <= 3'b000;
      // memory_array[27917] <= 3'b111;
      // memory_array[27918] <= 3'b000;
      // memory_array[27919] <= 3'b000;
      // memory_array[27920] <= 3'b000;
      // memory_array[27921] <= 3'b000;
      // memory_array[27922] <= 3'b101;
      // memory_array[27923] <= 3'b101;
      // memory_array[27924] <= 3'b000;
      // memory_array[27925] <= 3'b000;
      // memory_array[27926] <= 3'b111;
      // memory_array[27927] <= 3'b000;
      // memory_array[27928] <= 3'b101;
      // memory_array[27929] <= 3'b101;
      // memory_array[27930] <= 3'b000;
      // memory_array[27931] <= 3'b101;
      // memory_array[27932] <= 3'b000;
      // memory_array[27933] <= 3'b000;
      // memory_array[27934] <= 3'b111;
      // memory_array[27935] <= 3'b111;
      // memory_array[27936] <= 3'b101;
      // memory_array[27937] <= 3'b000;
      // memory_array[27938] <= 3'b111;
      // memory_array[27939] <= 3'b111;
      // memory_array[27940] <= 3'b000;
      // memory_array[27941] <= 3'b000;
      // memory_array[27942] <= 3'b000;
      // memory_array[27943] <= 3'b000;
      // memory_array[27944] <= 3'b101;
      // memory_array[27945] <= 3'b101;
      // memory_array[27946] <= 3'b000;
      // memory_array[27947] <= 3'b000;
      // memory_array[27948] <= 3'b000;
      // memory_array[27949] <= 3'b000;
      // memory_array[27950] <= 3'b111;
      // memory_array[27951] <= 3'b000;
      // memory_array[27952] <= 3'b000;
      // memory_array[27953] <= 3'b101;
      // memory_array[27954] <= 3'b000;
      // memory_array[27955] <= 3'b000;
      // memory_array[27956] <= 3'b000;
      // memory_array[27957] <= 3'b000;
      // memory_array[27958] <= 3'b000;
      // memory_array[27959] <= 3'b101;
      // memory_array[27960] <= 3'b000;
      // memory_array[27961] <= 3'b000;
      // memory_array[27962] <= 3'b000;
      // memory_array[27963] <= 3'b111;
      // memory_array[27964] <= 3'b000;
      // memory_array[27965] <= 3'b000;
      // memory_array[27966] <= 3'b000;
      // memory_array[27967] <= 3'b000;
      // memory_array[27968] <= 3'b000;
      // memory_array[27969] <= 3'b101;
      // memory_array[27970] <= 3'b101;
      // memory_array[27971] <= 3'b000;
      // memory_array[27972] <= 3'b000;
      // memory_array[27973] <= 3'b101;
      // memory_array[27974] <= 3'b101;
      // memory_array[27975] <= 3'b000;
      // memory_array[27976] <= 3'b111;
      // memory_array[27977] <= 3'b000;
      // memory_array[27978] <= 3'b101;
      // memory_array[27979] <= 3'b111;
      // memory_array[27980] <= 3'b111;
      // memory_array[27981] <= 3'b101;
      // memory_array[27982] <= 3'b101;
      // memory_array[27983] <= 3'b000;
      // memory_array[27984] <= 3'b101;
      // memory_array[27985] <= 3'b101;
      // memory_array[27986] <= 3'b000;
      // memory_array[27987] <= 3'b000;
      // memory_array[27988] <= 3'b111;
      // memory_array[27989] <= 3'b101;
      // memory_array[27990] <= 3'b101;
      // memory_array[27991] <= 3'b101;
      // memory_array[27992] <= 3'b111;
      // memory_array[27993] <= 3'b111;
      // memory_array[27994] <= 3'b111;
      // memory_array[27995] <= 3'b101;
      // memory_array[27996] <= 3'b101;
      // memory_array[27997] <= 3'b111;
      // memory_array[27998] <= 3'b111;
      // memory_array[27999] <= 3'b111;
      // memory_array[28000] <= 3'b111;
      // memory_array[28001] <= 3'b111;
      // memory_array[28002] <= 3'b101;
      // memory_array[28003] <= 3'b101;
      // memory_array[28004] <= 3'b111;
      // memory_array[28005] <= 3'b111;
      // memory_array[28006] <= 3'b111;
      // memory_array[28007] <= 3'b111;
      // memory_array[28008] <= 3'b101;
      // memory_array[28009] <= 3'b101;
      // memory_array[28010] <= 3'b000;
      // memory_array[28011] <= 3'b101;
      // memory_array[28012] <= 3'b000;
      // memory_array[28013] <= 3'b101;
      // memory_array[28014] <= 3'b111;
      // memory_array[28015] <= 3'b111;
      // memory_array[28016] <= 3'b101;
      // memory_array[28017] <= 3'b101;
      // memory_array[28018] <= 3'b000;
      // memory_array[28019] <= 3'b101;
      // memory_array[28020] <= 3'b101;
      // memory_array[28021] <= 3'b000;
      // memory_array[28022] <= 3'b000;
      // memory_array[28023] <= 3'b111;
      // memory_array[28024] <= 3'b101;
      // memory_array[28025] <= 3'b101;
      // memory_array[28026] <= 3'b101;
      // memory_array[28027] <= 3'b000;
      // memory_array[28028] <= 3'b000;
      // memory_array[28029] <= 3'b000;
      // memory_array[28030] <= 3'b101;
      // memory_array[28031] <= 3'b111;
      // memory_array[28032] <= 3'b000;
      // memory_array[28033] <= 3'b000;
      // memory_array[28034] <= 3'b111;
      // memory_array[28035] <= 3'b111;
      // memory_array[28036] <= 3'b101;
      // memory_array[28037] <= 3'b000;
      // memory_array[28038] <= 3'b111;
      // memory_array[28039] <= 3'b000;
      // memory_array[28040] <= 3'b000;
      // memory_array[28041] <= 3'b000;
      // memory_array[28042] <= 3'b000;
      // memory_array[28043] <= 3'b000;
      // memory_array[28044] <= 3'b000;
      // memory_array[28045] <= 3'b101;
      // memory_array[28046] <= 3'b000;
      // memory_array[28047] <= 3'b000;
      // memory_array[28048] <= 3'b000;
      // memory_array[28049] <= 3'b000;
      // memory_array[28050] <= 3'b101;
      // memory_array[28051] <= 3'b000;
      // memory_array[28052] <= 3'b000;
      // memory_array[28053] <= 3'b000;
      // memory_array[28054] <= 3'b000;
      // memory_array[28055] <= 3'b000;
      // memory_array[28056] <= 3'b000;
      // memory_array[28057] <= 3'b000;
      // memory_array[28058] <= 3'b000;
      // memory_array[28059] <= 3'b111;
      // memory_array[28060] <= 3'b000;
      // memory_array[28061] <= 3'b000;
      // memory_array[28062] <= 3'b000;
      // memory_array[28063] <= 3'b000;
      // memory_array[28064] <= 3'b000;
      // memory_array[28065] <= 3'b101;
      // memory_array[28066] <= 3'b000;
      // memory_array[28067] <= 3'b000;
      // memory_array[28068] <= 3'b111;
      // memory_array[28069] <= 3'b000;
      // memory_array[28070] <= 3'b000;
      // memory_array[28071] <= 3'b111;
      // memory_array[28072] <= 3'b000;
      // memory_array[28073] <= 3'b000;
      // memory_array[28074] <= 3'b000;
      // memory_array[28075] <= 3'b000;
      // memory_array[28076] <= 3'b111;
      // memory_array[28077] <= 3'b000;
      // memory_array[28078] <= 3'b000;
      // memory_array[28079] <= 3'b101;
      // memory_array[28080] <= 3'b111;
      // memory_array[28081] <= 3'b000;
      // memory_array[28082] <= 3'b111;
      // memory_array[28083] <= 3'b111;
      // memory_array[28084] <= 3'b000;
      // memory_array[28085] <= 3'b111;
      // memory_array[28086] <= 3'b000;
      // memory_array[28087] <= 3'b111;
      // memory_array[28088] <= 3'b111;
      // memory_array[28089] <= 3'b111;
      // memory_array[28090] <= 3'b111;
      // memory_array[28091] <= 3'b000;
      // memory_array[28092] <= 3'b111;
      // memory_array[28093] <= 3'b000;
      // memory_array[28094] <= 3'b111;
      // memory_array[28095] <= 3'b000;
      // memory_array[28096] <= 3'b111;
      // memory_array[28097] <= 3'b000;
      // memory_array[28098] <= 3'b101;
      // memory_array[28099] <= 3'b101;
      // memory_array[28100] <= 3'b101;
      // memory_array[28101] <= 3'b000;
      // memory_array[28102] <= 3'b111;
      // memory_array[28103] <= 3'b000;
      // memory_array[28104] <= 3'b000;
      // memory_array[28105] <= 3'b000;
      // memory_array[28106] <= 3'b000;
      // memory_array[28107] <= 3'b101;
      // memory_array[28108] <= 3'b000;
      // memory_array[28109] <= 3'b000;
      // memory_array[28110] <= 3'b000;
      // memory_array[28111] <= 3'b000;
      // memory_array[28112] <= 3'b000;
      // memory_array[28113] <= 3'b000;
      // memory_array[28114] <= 3'b101;
      // memory_array[28115] <= 3'b000;
      // memory_array[28116] <= 3'b000;
      // memory_array[28117] <= 3'b111;
      // memory_array[28118] <= 3'b000;
      // memory_array[28119] <= 3'b000;
      // memory_array[28120] <= 3'b000;
      // memory_array[28121] <= 3'b000;
      // memory_array[28122] <= 3'b101;
      // memory_array[28123] <= 3'b101;
      // memory_array[28124] <= 3'b000;
      // memory_array[28125] <= 3'b000;
      // memory_array[28126] <= 3'b111;
      // memory_array[28127] <= 3'b000;
      // memory_array[28128] <= 3'b101;
      // memory_array[28129] <= 3'b101;
      // memory_array[28130] <= 3'b000;
      // memory_array[28131] <= 3'b101;
      // memory_array[28132] <= 3'b000;
      // memory_array[28133] <= 3'b000;
      // memory_array[28134] <= 3'b111;
      // memory_array[28135] <= 3'b111;
      // memory_array[28136] <= 3'b101;
      // memory_array[28137] <= 3'b000;
      // memory_array[28138] <= 3'b111;
      // memory_array[28139] <= 3'b111;
      // memory_array[28140] <= 3'b000;
      // memory_array[28141] <= 3'b000;
      // memory_array[28142] <= 3'b000;
      // memory_array[28143] <= 3'b000;
      // memory_array[28144] <= 3'b101;
      // memory_array[28145] <= 3'b101;
      // memory_array[28146] <= 3'b000;
      // memory_array[28147] <= 3'b000;
      // memory_array[28148] <= 3'b000;
      // memory_array[28149] <= 3'b000;
      // memory_array[28150] <= 3'b111;
      // memory_array[28151] <= 3'b000;
      // memory_array[28152] <= 3'b000;
      // memory_array[28153] <= 3'b101;
      // memory_array[28154] <= 3'b000;
      // memory_array[28155] <= 3'b000;
      // memory_array[28156] <= 3'b000;
      // memory_array[28157] <= 3'b000;
      // memory_array[28158] <= 3'b000;
      // memory_array[28159] <= 3'b101;
      // memory_array[28160] <= 3'b000;
      // memory_array[28161] <= 3'b000;
      // memory_array[28162] <= 3'b000;
      // memory_array[28163] <= 3'b111;
      // memory_array[28164] <= 3'b000;
      // memory_array[28165] <= 3'b000;
      // memory_array[28166] <= 3'b000;
      // memory_array[28167] <= 3'b000;
      // memory_array[28168] <= 3'b000;
      // memory_array[28169] <= 3'b101;
      // memory_array[28170] <= 3'b101;
      // memory_array[28171] <= 3'b000;
      // memory_array[28172] <= 3'b000;
      // memory_array[28173] <= 3'b101;
      // memory_array[28174] <= 3'b101;
      // memory_array[28175] <= 3'b000;
      // memory_array[28176] <= 3'b111;
      // memory_array[28177] <= 3'b000;
      // memory_array[28178] <= 3'b101;
      // memory_array[28179] <= 3'b111;
      // memory_array[28180] <= 3'b111;
      // memory_array[28181] <= 3'b101;
      // memory_array[28182] <= 3'b101;
      // memory_array[28183] <= 3'b000;
      // memory_array[28184] <= 3'b101;
      // memory_array[28185] <= 3'b101;
      // memory_array[28186] <= 3'b000;
      // memory_array[28187] <= 3'b000;
      // memory_array[28188] <= 3'b111;
      // memory_array[28189] <= 3'b101;
      // memory_array[28190] <= 3'b101;
      // memory_array[28191] <= 3'b101;
      // memory_array[28192] <= 3'b111;
      // memory_array[28193] <= 3'b111;
      // memory_array[28194] <= 3'b111;
      // memory_array[28195] <= 3'b101;
      // memory_array[28196] <= 3'b101;
      // memory_array[28197] <= 3'b111;
      // memory_array[28198] <= 3'b111;
      // memory_array[28199] <= 3'b111;
      // memory_array[28200] <= 3'b111;
      // memory_array[28201] <= 3'b111;
      // memory_array[28202] <= 3'b101;
      // memory_array[28203] <= 3'b101;
      // memory_array[28204] <= 3'b111;
      // memory_array[28205] <= 3'b111;
      // memory_array[28206] <= 3'b111;
      // memory_array[28207] <= 3'b111;
      // memory_array[28208] <= 3'b101;
      // memory_array[28209] <= 3'b101;
      // memory_array[28210] <= 3'b000;
      // memory_array[28211] <= 3'b000;
      // memory_array[28212] <= 3'b101;
      // memory_array[28213] <= 3'b111;
      // memory_array[28214] <= 3'b111;
      // memory_array[28215] <= 3'b101;
      // memory_array[28216] <= 3'b000;
      // memory_array[28217] <= 3'b111;
      // memory_array[28218] <= 3'b111;
      // memory_array[28219] <= 3'b101;
      // memory_array[28220] <= 3'b000;
      // memory_array[28221] <= 3'b101;
      // memory_array[28222] <= 3'b111;
      // memory_array[28223] <= 3'b111;
      // memory_array[28224] <= 3'b101;
      // memory_array[28225] <= 3'b101;
      // memory_array[28226] <= 3'b101;
      // memory_array[28227] <= 3'b101;
      // memory_array[28228] <= 3'b101;
      // memory_array[28229] <= 3'b101;
      // memory_array[28230] <= 3'b000;
      // memory_array[28231] <= 3'b111;
      // memory_array[28232] <= 3'b111;
      // memory_array[28233] <= 3'b111;
      // memory_array[28234] <= 3'b000;
      // memory_array[28235] <= 3'b111;
      // memory_array[28236] <= 3'b000;
      // memory_array[28237] <= 3'b111;
      // memory_array[28238] <= 3'b111;
      // memory_array[28239] <= 3'b111;
      // memory_array[28240] <= 3'b111;
      // memory_array[28241] <= 3'b000;
      // memory_array[28242] <= 3'b111;
      // memory_array[28243] <= 3'b000;
      // memory_array[28244] <= 3'b111;
      // memory_array[28245] <= 3'b111;
      // memory_array[28246] <= 3'b000;
      // memory_array[28247] <= 3'b111;
      // memory_array[28248] <= 3'b000;
      // memory_array[28249] <= 3'b111;
      // memory_array[28250] <= 3'b111;
      // memory_array[28251] <= 3'b000;
      // memory_array[28252] <= 3'b111;
      // memory_array[28253] <= 3'b000;
      // memory_array[28254] <= 3'b000;
      // memory_array[28255] <= 3'b111;
      // memory_array[28256] <= 3'b000;
      // memory_array[28257] <= 3'b000;
      // memory_array[28258] <= 3'b111;
      // memory_array[28259] <= 3'b111;
      // memory_array[28260] <= 3'b000;
      // memory_array[28261] <= 3'b111;
      // memory_array[28262] <= 3'b000;
      // memory_array[28263] <= 3'b111;
      // memory_array[28264] <= 3'b000;
      // memory_array[28265] <= 3'b000;
      // memory_array[28266] <= 3'b111;
      // memory_array[28267] <= 3'b000;
      // memory_array[28268] <= 3'b111;
      // memory_array[28269] <= 3'b000;
      // memory_array[28270] <= 3'b000;
      // memory_array[28271] <= 3'b111;
      // memory_array[28272] <= 3'b000;
      // memory_array[28273] <= 3'b111;
      // memory_array[28274] <= 3'b000;
      // memory_array[28275] <= 3'b000;
      // memory_array[28276] <= 3'b111;
      // memory_array[28277] <= 3'b000;
      // memory_array[28278] <= 3'b000;
      // memory_array[28279] <= 3'b000;
      // memory_array[28280] <= 3'b101;
      // memory_array[28281] <= 3'b101;
      // memory_array[28282] <= 3'b111;
      // memory_array[28283] <= 3'b111;
      // memory_array[28284] <= 3'b101;
      // memory_array[28285] <= 3'b000;
      // memory_array[28286] <= 3'b111;
      // memory_array[28287] <= 3'b111;
      // memory_array[28288] <= 3'b111;
      // memory_array[28289] <= 3'b000;
      // memory_array[28290] <= 3'b111;
      // memory_array[28291] <= 3'b111;
      // memory_array[28292] <= 3'b111;
      // memory_array[28293] <= 3'b000;
      // memory_array[28294] <= 3'b111;
      // memory_array[28295] <= 3'b000;
      // memory_array[28296] <= 3'b111;
      // memory_array[28297] <= 3'b000;
      // memory_array[28298] <= 3'b101;
      // memory_array[28299] <= 3'b101;
      // memory_array[28300] <= 3'b101;
      // memory_array[28301] <= 3'b000;
      // memory_array[28302] <= 3'b111;
      // memory_array[28303] <= 3'b000;
      // memory_array[28304] <= 3'b111;
      // memory_array[28305] <= 3'b111;
      // memory_array[28306] <= 3'b000;
      // memory_array[28307] <= 3'b111;
      // memory_array[28308] <= 3'b000;
      // memory_array[28309] <= 3'b111;
      // memory_array[28310] <= 3'b111;
      // memory_array[28311] <= 3'b000;
      // memory_array[28312] <= 3'b111;
      // memory_array[28313] <= 3'b000;
      // memory_array[28314] <= 3'b111;
      // memory_array[28315] <= 3'b000;
      // memory_array[28316] <= 3'b111;
      // memory_array[28317] <= 3'b111;
      // memory_array[28318] <= 3'b000;
      // memory_array[28319] <= 3'b000;
      // memory_array[28320] <= 3'b000;
      // memory_array[28321] <= 3'b000;
      // memory_array[28322] <= 3'b111;
      // memory_array[28323] <= 3'b000;
      // memory_array[28324] <= 3'b000;
      // memory_array[28325] <= 3'b111;
      // memory_array[28326] <= 3'b111;
      // memory_array[28327] <= 3'b111;
      // memory_array[28328] <= 3'b111;
      // memory_array[28329] <= 3'b101;
      // memory_array[28330] <= 3'b000;
      // memory_array[28331] <= 3'b000;
      // memory_array[28332] <= 3'b101;
      // memory_array[28333] <= 3'b000;
      // memory_array[28334] <= 3'b000;
      // memory_array[28335] <= 3'b111;
      // memory_array[28336] <= 3'b000;
      // memory_array[28337] <= 3'b111;
      // memory_array[28338] <= 3'b000;
      // memory_array[28339] <= 3'b111;
      // memory_array[28340] <= 3'b000;
      // memory_array[28341] <= 3'b111;
      // memory_array[28342] <= 3'b000;
      // memory_array[28343] <= 3'b000;
      // memory_array[28344] <= 3'b000;
      // memory_array[28345] <= 3'b000;
      // memory_array[28346] <= 3'b111;
      // memory_array[28347] <= 3'b000;
      // memory_array[28348] <= 3'b111;
      // memory_array[28349] <= 3'b000;
      // memory_array[28350] <= 3'b111;
      // memory_array[28351] <= 3'b111;
      // memory_array[28352] <= 3'b111;
      // memory_array[28353] <= 3'b111;
      // memory_array[28354] <= 3'b000;
      // memory_array[28355] <= 3'b000;
      // memory_array[28356] <= 3'b111;
      // memory_array[28357] <= 3'b000;
      // memory_array[28358] <= 3'b111;
      // memory_array[28359] <= 3'b000;
      // memory_array[28360] <= 3'b000;
      // memory_array[28361] <= 3'b111;
      // memory_array[28362] <= 3'b000;
      // memory_array[28363] <= 3'b111;
      // memory_array[28364] <= 3'b000;
      // memory_array[28365] <= 3'b000;
      // memory_array[28366] <= 3'b111;
      // memory_array[28367] <= 3'b000;
      // memory_array[28368] <= 3'b111;
      // memory_array[28369] <= 3'b000;
      // memory_array[28370] <= 3'b101;
      // memory_array[28371] <= 3'b101;
      // memory_array[28372] <= 3'b000;
      // memory_array[28373] <= 3'b101;
      // memory_array[28374] <= 3'b101;
      // memory_array[28375] <= 3'b000;
      // memory_array[28376] <= 3'b000;
      // memory_array[28377] <= 3'b101;
      // memory_array[28378] <= 3'b111;
      // memory_array[28379] <= 3'b111;
      // memory_array[28380] <= 3'b101;
      // memory_array[28381] <= 3'b000;
      // memory_array[28382] <= 3'b111;
      // memory_array[28383] <= 3'b111;
      // memory_array[28384] <= 3'b101;
      // memory_array[28385] <= 3'b000;
      // memory_array[28386] <= 3'b101;
      // memory_array[28387] <= 3'b111;
      // memory_array[28388] <= 3'b111;
      // memory_array[28389] <= 3'b101;
      // memory_array[28390] <= 3'b101;
      // memory_array[28391] <= 3'b101;
      // memory_array[28392] <= 3'b111;
      // memory_array[28393] <= 3'b101;
      // memory_array[28394] <= 3'b101;
      // memory_array[28395] <= 3'b111;
      // memory_array[28396] <= 3'b111;
      // memory_array[28397] <= 3'b101;
      // memory_array[28398] <= 3'b101;
      // memory_array[28399] <= 3'b111;
      // memory_array[28400] <= 3'b111;
      // memory_array[28401] <= 3'b111;
      // memory_array[28402] <= 3'b101;
      // memory_array[28403] <= 3'b101;
      // memory_array[28404] <= 3'b111;
      // memory_array[28405] <= 3'b101;
      // memory_array[28406] <= 3'b111;
      // memory_array[28407] <= 3'b111;
      // memory_array[28408] <= 3'b101;
      // memory_array[28409] <= 3'b101;
      // memory_array[28410] <= 3'b000;
      // memory_array[28411] <= 3'b000;
      // memory_array[28412] <= 3'b000;
      // memory_array[28413] <= 3'b101;
      // memory_array[28414] <= 3'b000;
      // memory_array[28415] <= 3'b101;
      // memory_array[28416] <= 3'b101;
      // memory_array[28417] <= 3'b101;
      // memory_array[28418] <= 3'b000;
      // memory_array[28419] <= 3'b101;
      // memory_array[28420] <= 3'b000;
      // memory_array[28421] <= 3'b000;
      // memory_array[28422] <= 3'b101;
      // memory_array[28423] <= 3'b111;
      // memory_array[28424] <= 3'b101;
      // memory_array[28425] <= 3'b101;
      // memory_array[28426] <= 3'b101;
      // memory_array[28427] <= 3'b000;
      // memory_array[28428] <= 3'b000;
      // memory_array[28429] <= 3'b000;
      // memory_array[28430] <= 3'b000;
      // memory_array[28431] <= 3'b111;
      // memory_array[28432] <= 3'b000;
      // memory_array[28433] <= 3'b000;
      // memory_array[28434] <= 3'b111;
      // memory_array[28435] <= 3'b111;
      // memory_array[28436] <= 3'b101;
      // memory_array[28437] <= 3'b000;
      // memory_array[28438] <= 3'b111;
      // memory_array[28439] <= 3'b000;
      // memory_array[28440] <= 3'b000;
      // memory_array[28441] <= 3'b000;
      // memory_array[28442] <= 3'b111;
      // memory_array[28443] <= 3'b000;
      // memory_array[28444] <= 3'b111;
      // memory_array[28445] <= 3'b111;
      // memory_array[28446] <= 3'b000;
      // memory_array[28447] <= 3'b111;
      // memory_array[28448] <= 3'b000;
      // memory_array[28449] <= 3'b111;
      // memory_array[28450] <= 3'b000;
      // memory_array[28451] <= 3'b111;
      // memory_array[28452] <= 3'b111;
      // memory_array[28453] <= 3'b111;
      // memory_array[28454] <= 3'b111;
      // memory_array[28455] <= 3'b111;
      // memory_array[28456] <= 3'b000;
      // memory_array[28457] <= 3'b000;
      // memory_array[28458] <= 3'b111;
      // memory_array[28459] <= 3'b000;
      // memory_array[28460] <= 3'b000;
      // memory_array[28461] <= 3'b101;
      // memory_array[28462] <= 3'b000;
      // memory_array[28463] <= 3'b111;
      // memory_array[28464] <= 3'b000;
      // memory_array[28465] <= 3'b000;
      // memory_array[28466] <= 3'b111;
      // memory_array[28467] <= 3'b111;
      // memory_array[28468] <= 3'b111;
      // memory_array[28469] <= 3'b000;
      // memory_array[28470] <= 3'b000;
      // memory_array[28471] <= 3'b111;
      // memory_array[28472] <= 3'b000;
      // memory_array[28473] <= 3'b111;
      // memory_array[28474] <= 3'b000;
      // memory_array[28475] <= 3'b000;
      // memory_array[28476] <= 3'b111;
      // memory_array[28477] <= 3'b111;
      // memory_array[28478] <= 3'b111;
      // memory_array[28479] <= 3'b101;
      // memory_array[28480] <= 3'b101;
      // memory_array[28481] <= 3'b000;
      // memory_array[28482] <= 3'b111;
      // memory_array[28483] <= 3'b111;
      // memory_array[28484] <= 3'b000;
      // memory_array[28485] <= 3'b000;
      // memory_array[28486] <= 3'b111;
      // memory_array[28487] <= 3'b000;
      // memory_array[28488] <= 3'b101;
      // memory_array[28489] <= 3'b000;
      // memory_array[28490] <= 3'b000;
      // memory_array[28491] <= 3'b111;
      // memory_array[28492] <= 3'b101;
      // memory_array[28493] <= 3'b000;
      // memory_array[28494] <= 3'b111;
      // memory_array[28495] <= 3'b000;
      // memory_array[28496] <= 3'b111;
      // memory_array[28497] <= 3'b000;
      // memory_array[28498] <= 3'b101;
      // memory_array[28499] <= 3'b101;
      // memory_array[28500] <= 3'b101;
      // memory_array[28501] <= 3'b000;
      // memory_array[28502] <= 3'b111;
      // memory_array[28503] <= 3'b000;
      // memory_array[28504] <= 3'b111;
      // memory_array[28505] <= 3'b111;
      // memory_array[28506] <= 3'b000;
      // memory_array[28507] <= 3'b111;
      // memory_array[28508] <= 3'b000;
      // memory_array[28509] <= 3'b111;
      // memory_array[28510] <= 3'b111;
      // memory_array[28511] <= 3'b000;
      // memory_array[28512] <= 3'b000;
      // memory_array[28513] <= 3'b000;
      // memory_array[28514] <= 3'b111;
      // memory_array[28515] <= 3'b000;
      // memory_array[28516] <= 3'b111;
      // memory_array[28517] <= 3'b111;
      // memory_array[28518] <= 3'b000;
      // memory_array[28519] <= 3'b111;
      // memory_array[28520] <= 3'b111;
      // memory_array[28521] <= 3'b000;
      // memory_array[28522] <= 3'b111;
      // memory_array[28523] <= 3'b000;
      // memory_array[28524] <= 3'b000;
      // memory_array[28525] <= 3'b111;
      // memory_array[28526] <= 3'b000;
      // memory_array[28527] <= 3'b111;
      // memory_array[28528] <= 3'b111;
      // memory_array[28529] <= 3'b000;
      // memory_array[28530] <= 3'b000;
      // memory_array[28531] <= 3'b000;
      // memory_array[28532] <= 3'b000;
      // memory_array[28533] <= 3'b000;
      // memory_array[28534] <= 3'b000;
      // memory_array[28535] <= 3'b000;
      // memory_array[28536] <= 3'b111;
      // memory_array[28537] <= 3'b000;
      // memory_array[28538] <= 3'b000;
      // memory_array[28539] <= 3'b111;
      // memory_array[28540] <= 3'b000;
      // memory_array[28541] <= 3'b111;
      // memory_array[28542] <= 3'b000;
      // memory_array[28543] <= 3'b000;
      // memory_array[28544] <= 3'b000;
      // memory_array[28545] <= 3'b000;
      // memory_array[28546] <= 3'b111;
      // memory_array[28547] <= 3'b000;
      // memory_array[28548] <= 3'b000;
      // memory_array[28549] <= 3'b000;
      // memory_array[28550] <= 3'b111;
      // memory_array[28551] <= 3'b000;
      // memory_array[28552] <= 3'b111;
      // memory_array[28553] <= 3'b111;
      // memory_array[28554] <= 3'b000;
      // memory_array[28555] <= 3'b000;
      // memory_array[28556] <= 3'b111;
      // memory_array[28557] <= 3'b000;
      // memory_array[28558] <= 3'b111;
      // memory_array[28559] <= 3'b000;
      // memory_array[28560] <= 3'b000;
      // memory_array[28561] <= 3'b111;
      // memory_array[28562] <= 3'b000;
      // memory_array[28563] <= 3'b000;
      // memory_array[28564] <= 3'b000;
      // memory_array[28565] <= 3'b000;
      // memory_array[28566] <= 3'b111;
      // memory_array[28567] <= 3'b000;
      // memory_array[28568] <= 3'b101;
      // memory_array[28569] <= 3'b101;
      // memory_array[28570] <= 3'b000;
      // memory_array[28571] <= 3'b000;
      // memory_array[28572] <= 3'b000;
      // memory_array[28573] <= 3'b000;
      // memory_array[28574] <= 3'b101;
      // memory_array[28575] <= 3'b000;
      // memory_array[28576] <= 3'b000;
      // memory_array[28577] <= 3'b000;
      // memory_array[28578] <= 3'b101;
      // memory_array[28579] <= 3'b000;
      // memory_array[28580] <= 3'b101;
      // memory_array[28581] <= 3'b101;
      // memory_array[28582] <= 3'b101;
      // memory_array[28583] <= 3'b000;
      // memory_array[28584] <= 3'b101;
      // memory_array[28585] <= 3'b000;
      // memory_array[28586] <= 3'b000;
      // memory_array[28587] <= 3'b101;
      // memory_array[28588] <= 3'b111;
      // memory_array[28589] <= 3'b101;
      // memory_array[28590] <= 3'b101;
      // memory_array[28591] <= 3'b101;
      // memory_array[28592] <= 3'b111;
      // memory_array[28593] <= 3'b111;
      // memory_array[28594] <= 3'b111;
      // memory_array[28595] <= 3'b101;
      // memory_array[28596] <= 3'b101;
      // memory_array[28597] <= 3'b111;
      // memory_array[28598] <= 3'b111;
      // memory_array[28599] <= 3'b111;
      // memory_array[28600] <= 3'b111;
      // memory_array[28601] <= 3'b111;
      // memory_array[28602] <= 3'b101;
      // memory_array[28603] <= 3'b101;
      // memory_array[28604] <= 3'b101;
      // memory_array[28605] <= 3'b101;
      // memory_array[28606] <= 3'b111;
      // memory_array[28607] <= 3'b111;
      // memory_array[28608] <= 3'b101;
      // memory_array[28609] <= 3'b101;
      // memory_array[28610] <= 3'b000;
      // memory_array[28611] <= 3'b000;
      // memory_array[28612] <= 3'b101;
      // memory_array[28613] <= 3'b000;
      // memory_array[28614] <= 3'b111;
      // memory_array[28615] <= 3'b101;
      // memory_array[28616] <= 3'b101;
      // memory_array[28617] <= 3'b111;
      // memory_array[28618] <= 3'b101;
      // memory_array[28619] <= 3'b111;
      // memory_array[28620] <= 3'b101;
      // memory_array[28621] <= 3'b000;
      // memory_array[28622] <= 3'b111;
      // memory_array[28623] <= 3'b101;
      // memory_array[28624] <= 3'b111;
      // memory_array[28625] <= 3'b101;
      // memory_array[28626] <= 3'b101;
      // memory_array[28627] <= 3'b101;
      // memory_array[28628] <= 3'b101;
      // memory_array[28629] <= 3'b101;
      // memory_array[28630] <= 3'b000;
      // memory_array[28631] <= 3'b000;
      // memory_array[28632] <= 3'b111;
      // memory_array[28633] <= 3'b111;
      // memory_array[28634] <= 3'b111;
      // memory_array[28635] <= 3'b000;
      // memory_array[28636] <= 3'b000;
      // memory_array[28637] <= 3'b000;
      // memory_array[28638] <= 3'b000;
      // memory_array[28639] <= 3'b111;
      // memory_array[28640] <= 3'b111;
      // memory_array[28641] <= 3'b000;
      // memory_array[28642] <= 3'b111;
      // memory_array[28643] <= 3'b111;
      // memory_array[28644] <= 3'b111;
      // memory_array[28645] <= 3'b000;
      // memory_array[28646] <= 3'b000;
      // memory_array[28647] <= 3'b111;
      // memory_array[28648] <= 3'b111;
      // memory_array[28649] <= 3'b000;
      // memory_array[28650] <= 3'b000;
      // memory_array[28651] <= 3'b101;
      // memory_array[28652] <= 3'b000;
      // memory_array[28653] <= 3'b111;
      // memory_array[28654] <= 3'b111;
      // memory_array[28655] <= 3'b000;
      // memory_array[28656] <= 3'b000;
      // memory_array[28657] <= 3'b111;
      // memory_array[28658] <= 3'b111;
      // memory_array[28659] <= 3'b111;
      // memory_array[28660] <= 3'b000;
      // memory_array[28661] <= 3'b101;
      // memory_array[28662] <= 3'b111;
      // memory_array[28663] <= 3'b111;
      // memory_array[28664] <= 3'b111;
      // memory_array[28665] <= 3'b000;
      // memory_array[28666] <= 3'b111;
      // memory_array[28667] <= 3'b000;
      // memory_array[28668] <= 3'b111;
      // memory_array[28669] <= 3'b000;
      // memory_array[28670] <= 3'b111;
      // memory_array[28671] <= 3'b111;
      // memory_array[28672] <= 3'b000;
      // memory_array[28673] <= 3'b111;
      // memory_array[28674] <= 3'b111;
      // memory_array[28675] <= 3'b000;
      // memory_array[28676] <= 3'b111;
      // memory_array[28677] <= 3'b111;
      // memory_array[28678] <= 3'b000;
      // memory_array[28679] <= 3'b000;
      // memory_array[28680] <= 3'b000;
      // memory_array[28681] <= 3'b000;
      // memory_array[28682] <= 3'b111;
      // memory_array[28683] <= 3'b111;
      // memory_array[28684] <= 3'b000;
      // memory_array[28685] <= 3'b000;
      // memory_array[28686] <= 3'b111;
      // memory_array[28687] <= 3'b111;
      // memory_array[28688] <= 3'b111;
      // memory_array[28689] <= 3'b000;
      // memory_array[28690] <= 3'b111;
      // memory_array[28691] <= 3'b000;
      // memory_array[28692] <= 3'b101;
      // memory_array[28693] <= 3'b101;
      // memory_array[28694] <= 3'b111;
      // memory_array[28695] <= 3'b111;
      // memory_array[28696] <= 3'b111;
      // memory_array[28697] <= 3'b000;
      // memory_array[28698] <= 3'b101;
      // memory_array[28699] <= 3'b101;
      // memory_array[28700] <= 3'b101;
      // memory_array[28701] <= 3'b000;
      // memory_array[28702] <= 3'b111;
      // memory_array[28703] <= 3'b000;
      // memory_array[28704] <= 3'b000;
      // memory_array[28705] <= 3'b111;
      // memory_array[28706] <= 3'b111;
      // memory_array[28707] <= 3'b000;
      // memory_array[28708] <= 3'b000;
      // memory_array[28709] <= 3'b111;
      // memory_array[28710] <= 3'b111;
      // memory_array[28711] <= 3'b000;
      // memory_array[28712] <= 3'b000;
      // memory_array[28713] <= 3'b000;
      // memory_array[28714] <= 3'b111;
      // memory_array[28715] <= 3'b111;
      // memory_array[28716] <= 3'b000;
      // memory_array[28717] <= 3'b111;
      // memory_array[28718] <= 3'b111;
      // memory_array[28719] <= 3'b000;
      // memory_array[28720] <= 3'b111;
      // memory_array[28721] <= 3'b111;
      // memory_array[28722] <= 3'b111;
      // memory_array[28723] <= 3'b111;
      // memory_array[28724] <= 3'b111;
      // memory_array[28725] <= 3'b111;
      // memory_array[28726] <= 3'b111;
      // memory_array[28727] <= 3'b111;
      // memory_array[28728] <= 3'b111;
      // memory_array[28729] <= 3'b000;
      // memory_array[28730] <= 3'b000;
      // memory_array[28731] <= 3'b000;
      // memory_array[28732] <= 3'b000;
      // memory_array[28733] <= 3'b111;
      // memory_array[28734] <= 3'b111;
      // memory_array[28735] <= 3'b000;
      // memory_array[28736] <= 3'b111;
      // memory_array[28737] <= 3'b000;
      // memory_array[28738] <= 3'b111;
      // memory_array[28739] <= 3'b111;
      // memory_array[28740] <= 3'b111;
      // memory_array[28741] <= 3'b000;
      // memory_array[28742] <= 3'b111;
      // memory_array[28743] <= 3'b111;
      // memory_array[28744] <= 3'b000;
      // memory_array[28745] <= 3'b101;
      // memory_array[28746] <= 3'b111;
      // memory_array[28747] <= 3'b111;
      // memory_array[28748] <= 3'b111;
      // memory_array[28749] <= 3'b111;
      // memory_array[28750] <= 3'b111;
      // memory_array[28751] <= 3'b111;
      // memory_array[28752] <= 3'b111;
      // memory_array[28753] <= 3'b111;
      // memory_array[28754] <= 3'b000;
      // memory_array[28755] <= 3'b111;
      // memory_array[28756] <= 3'b111;
      // memory_array[28757] <= 3'b000;
      // memory_array[28758] <= 3'b111;
      // memory_array[28759] <= 3'b111;
      // memory_array[28760] <= 3'b000;
      // memory_array[28761] <= 3'b111;
      // memory_array[28762] <= 3'b111;
      // memory_array[28763] <= 3'b111;
      // memory_array[28764] <= 3'b000;
      // memory_array[28765] <= 3'b111;
      // memory_array[28766] <= 3'b111;
      // memory_array[28767] <= 3'b000;
      // memory_array[28768] <= 3'b000;
      // memory_array[28769] <= 3'b101;
      // memory_array[28770] <= 3'b101;
      // memory_array[28771] <= 3'b101;
      // memory_array[28772] <= 3'b000;
      // memory_array[28773] <= 3'b000;
      // memory_array[28774] <= 3'b101;
      // memory_array[28775] <= 3'b000;
      // memory_array[28776] <= 3'b000;
      // memory_array[28777] <= 3'b101;
      // memory_array[28778] <= 3'b000;
      // memory_array[28779] <= 3'b111;
      // memory_array[28780] <= 3'b101;
      // memory_array[28781] <= 3'b101;
      // memory_array[28782] <= 3'b111;
      // memory_array[28783] <= 3'b101;
      // memory_array[28784] <= 3'b111;
      // memory_array[28785] <= 3'b101;
      // memory_array[28786] <= 3'b000;
      // memory_array[28787] <= 3'b111;
      // memory_array[28788] <= 3'b101;
      // memory_array[28789] <= 3'b111;
      // memory_array[28790] <= 3'b101;
      // memory_array[28791] <= 3'b101;
      // memory_array[28792] <= 3'b111;
      // memory_array[28793] <= 3'b111;
      // memory_array[28794] <= 3'b111;
      // memory_array[28795] <= 3'b101;
      // memory_array[28796] <= 3'b101;
      // memory_array[28797] <= 3'b111;
      // memory_array[28798] <= 3'b111;
      // memory_array[28799] <= 3'b111;
      // memory_array[28800] <= 3'b111;
      // memory_array[28801] <= 3'b111;
      // memory_array[28802] <= 3'b101;
      // memory_array[28803] <= 3'b101;
      // memory_array[28804] <= 3'b111;
      // memory_array[28805] <= 3'b101;
      // memory_array[28806] <= 3'b111;
      // memory_array[28807] <= 3'b111;
      // memory_array[28808] <= 3'b101;
      // memory_array[28809] <= 3'b101;
      // memory_array[28810] <= 3'b000;
      // memory_array[28811] <= 3'b000;
      // memory_array[28812] <= 3'b000;
      // memory_array[28813] <= 3'b101;
      // memory_array[28814] <= 3'b101;
      // memory_array[28815] <= 3'b000;
      // memory_array[28816] <= 3'b101;
      // memory_array[28817] <= 3'b000;
      // memory_array[28818] <= 3'b000;
      // memory_array[28819] <= 3'b111;
      // memory_array[28820] <= 3'b000;
      // memory_array[28821] <= 3'b000;
      // memory_array[28822] <= 3'b101;
      // memory_array[28823] <= 3'b000;
      // memory_array[28824] <= 3'b101;
      // memory_array[28825] <= 3'b101;
      // memory_array[28826] <= 3'b101;
      // memory_array[28827] <= 3'b101;
      // memory_array[28828] <= 3'b101;
      // memory_array[28829] <= 3'b101;
      // memory_array[28830] <= 3'b101;
      // memory_array[28831] <= 3'b000;
      // memory_array[28832] <= 3'b000;
      // memory_array[28833] <= 3'b000;
      // memory_array[28834] <= 3'b000;
      // memory_array[28835] <= 3'b101;
      // memory_array[28836] <= 3'b000;
      // memory_array[28837] <= 3'b000;
      // memory_array[28838] <= 3'b000;
      // memory_array[28839] <= 3'b000;
      // memory_array[28840] <= 3'b000;
      // memory_array[28841] <= 3'b000;
      // memory_array[28842] <= 3'b000;
      // memory_array[28843] <= 3'b000;
      // memory_array[28844] <= 3'b000;
      // memory_array[28845] <= 3'b111;
      // memory_array[28846] <= 3'b000;
      // memory_array[28847] <= 3'b111;
      // memory_array[28848] <= 3'b000;
      // memory_array[28849] <= 3'b000;
      // memory_array[28850] <= 3'b000;
      // memory_array[28851] <= 3'b000;
      // memory_array[28852] <= 3'b000;
      // memory_array[28853] <= 3'b111;
      // memory_array[28854] <= 3'b000;
      // memory_array[28855] <= 3'b000;
      // memory_array[28856] <= 3'b101;
      // memory_array[28857] <= 3'b000;
      // memory_array[28858] <= 3'b000;
      // memory_array[28859] <= 3'b000;
      // memory_array[28860] <= 3'b000;
      // memory_array[28861] <= 3'b101;
      // memory_array[28862] <= 3'b000;
      // memory_array[28863] <= 3'b000;
      // memory_array[28864] <= 3'b000;
      // memory_array[28865] <= 3'b000;
      // memory_array[28866] <= 3'b111;
      // memory_array[28867] <= 3'b000;
      // memory_array[28868] <= 3'b111;
      // memory_array[28869] <= 3'b000;
      // memory_array[28870] <= 3'b000;
      // memory_array[28871] <= 3'b000;
      // memory_array[28872] <= 3'b000;
      // memory_array[28873] <= 3'b000;
      // memory_array[28874] <= 3'b000;
      // memory_array[28875] <= 3'b000;
      // memory_array[28876] <= 3'b000;
      // memory_array[28877] <= 3'b000;
      // memory_array[28878] <= 3'b000;
      // memory_array[28879] <= 3'b000;
      // memory_array[28880] <= 3'b000;
      // memory_array[28881] <= 3'b000;
      // memory_array[28882] <= 3'b000;
      // memory_array[28883] <= 3'b000;
      // memory_array[28884] <= 3'b000;
      // memory_array[28885] <= 3'b000;
      // memory_array[28886] <= 3'b000;
      // memory_array[28887] <= 3'b101;
      // memory_array[28888] <= 3'b101;
      // memory_array[28889] <= 3'b101;
      // memory_array[28890] <= 3'b000;
      // memory_array[28891] <= 3'b101;
      // memory_array[28892] <= 3'b101;
      // memory_array[28893] <= 3'b101;
      // memory_array[28894] <= 3'b000;
      // memory_array[28895] <= 3'b000;
      // memory_array[28896] <= 3'b000;
      // memory_array[28897] <= 3'b000;
      // memory_array[28898] <= 3'b101;
      // memory_array[28899] <= 3'b101;
      // memory_array[28900] <= 3'b101;
      // memory_array[28901] <= 3'b111;
      // memory_array[28902] <= 3'b000;
      // memory_array[28903] <= 3'b101;
      // memory_array[28904] <= 3'b101;
      // memory_array[28905] <= 3'b000;
      // memory_array[28906] <= 3'b000;
      // memory_array[28907] <= 3'b000;
      // memory_array[28908] <= 3'b000;
      // memory_array[28909] <= 3'b000;
      // memory_array[28910] <= 3'b000;
      // memory_array[28911] <= 3'b000;
      // memory_array[28912] <= 3'b000;
      // memory_array[28913] <= 3'b000;
      // memory_array[28914] <= 3'b000;
      // memory_array[28915] <= 3'b000;
      // memory_array[28916] <= 3'b101;
      // memory_array[28917] <= 3'b000;
      // memory_array[28918] <= 3'b000;
      // memory_array[28919] <= 3'b000;
      // memory_array[28920] <= 3'b000;
      // memory_array[28921] <= 3'b000;
      // memory_array[28922] <= 3'b000;
      // memory_array[28923] <= 3'b000;
      // memory_array[28924] <= 3'b000;
      // memory_array[28925] <= 3'b000;
      // memory_array[28926] <= 3'b000;
      // memory_array[28927] <= 3'b000;
      // memory_array[28928] <= 3'b000;
      // memory_array[28929] <= 3'b000;
      // memory_array[28930] <= 3'b000;
      // memory_array[28931] <= 3'b101;
      // memory_array[28932] <= 3'b000;
      // memory_array[28933] <= 3'b000;
      // memory_array[28934] <= 3'b000;
      // memory_array[28935] <= 3'b000;
      // memory_array[28936] <= 3'b000;
      // memory_array[28937] <= 3'b000;
      // memory_array[28938] <= 3'b000;
      // memory_array[28939] <= 3'b000;
      // memory_array[28940] <= 3'b000;
      // memory_array[28941] <= 3'b000;
      // memory_array[28942] <= 3'b000;
      // memory_array[28943] <= 3'b000;
      // memory_array[28944] <= 3'b000;
      // memory_array[28945] <= 3'b000;
      // memory_array[28946] <= 3'b000;
      // memory_array[28947] <= 3'b000;
      // memory_array[28948] <= 3'b000;
      // memory_array[28949] <= 3'b000;
      // memory_array[28950] <= 3'b000;
      // memory_array[28951] <= 3'b000;
      // memory_array[28952] <= 3'b000;
      // memory_array[28953] <= 3'b000;
      // memory_array[28954] <= 3'b000;
      // memory_array[28955] <= 3'b000;
      // memory_array[28956] <= 3'b000;
      // memory_array[28957] <= 3'b000;
      // memory_array[28958] <= 3'b000;
      // memory_array[28959] <= 3'b000;
      // memory_array[28960] <= 3'b000;
      // memory_array[28961] <= 3'b000;
      // memory_array[28962] <= 3'b000;
      // memory_array[28963] <= 3'b000;
      // memory_array[28964] <= 3'b000;
      // memory_array[28965] <= 3'b000;
      // memory_array[28966] <= 3'b000;
      // memory_array[28967] <= 3'b000;
      // memory_array[28968] <= 3'b101;
      // memory_array[28969] <= 3'b101;
      // memory_array[28970] <= 3'b101;
      // memory_array[28971] <= 3'b101;
      // memory_array[28972] <= 3'b000;
      // memory_array[28973] <= 3'b000;
      // memory_array[28974] <= 3'b101;
      // memory_array[28975] <= 3'b000;
      // memory_array[28976] <= 3'b101;
      // memory_array[28977] <= 3'b000;
      // memory_array[28978] <= 3'b101;
      // memory_array[28979] <= 3'b101;
      // memory_array[28980] <= 3'b000;
      // memory_array[28981] <= 3'b101;
      // memory_array[28982] <= 3'b000;
      // memory_array[28983] <= 3'b000;
      // memory_array[28984] <= 3'b111;
      // memory_array[28985] <= 3'b000;
      // memory_array[28986] <= 3'b000;
      // memory_array[28987] <= 3'b101;
      // memory_array[28988] <= 3'b000;
      // memory_array[28989] <= 3'b101;
      // memory_array[28990] <= 3'b101;
      // memory_array[28991] <= 3'b101;
      // memory_array[28992] <= 3'b111;
      // memory_array[28993] <= 3'b111;
      // memory_array[28994] <= 3'b111;
      // memory_array[28995] <= 3'b101;
      // memory_array[28996] <= 3'b101;
      // memory_array[28997] <= 3'b111;
      // memory_array[28998] <= 3'b111;
      // memory_array[28999] <= 3'b111;
      // memory_array[29000] <= 3'b111;
      // memory_array[29001] <= 3'b111;
      // memory_array[29002] <= 3'b101;
      // memory_array[29003] <= 3'b101;
      // memory_array[29004] <= 3'b111;
      // memory_array[29005] <= 3'b101;
      // memory_array[29006] <= 3'b111;
      // memory_array[29007] <= 3'b111;
      // memory_array[29008] <= 3'b101;
      // memory_array[29009] <= 3'b101;
      // memory_array[29010] <= 3'b101;
      // memory_array[29011] <= 3'b000;
      // memory_array[29012] <= 3'b000;
      // memory_array[29013] <= 3'b000;
      // memory_array[29014] <= 3'b101;
      // memory_array[29015] <= 3'b000;
      // memory_array[29016] <= 3'b101;
      // memory_array[29017] <= 3'b000;
      // memory_array[29018] <= 3'b000;
      // memory_array[29019] <= 3'b101;
      // memory_array[29020] <= 3'b000;
      // memory_array[29021] <= 3'b111;
      // memory_array[29022] <= 3'b101;
      // memory_array[29023] <= 3'b111;
      // memory_array[29024] <= 3'b101;
      // memory_array[29025] <= 3'b101;
      // memory_array[29026] <= 3'b101;
      // memory_array[29027] <= 3'b101;
      // memory_array[29028] <= 3'b101;
      // memory_array[29029] <= 3'b101;
      // memory_array[29030] <= 3'b101;
      // memory_array[29031] <= 3'b101;
      // memory_array[29032] <= 3'b101;
      // memory_array[29033] <= 3'b101;
      // memory_array[29034] <= 3'b101;
      // memory_array[29035] <= 3'b101;
      // memory_array[29036] <= 3'b101;
      // memory_array[29037] <= 3'b000;
      // memory_array[29038] <= 3'b000;
      // memory_array[29039] <= 3'b101;
      // memory_array[29040] <= 3'b101;
      // memory_array[29041] <= 3'b101;
      // memory_array[29042] <= 3'b101;
      // memory_array[29043] <= 3'b101;
      // memory_array[29044] <= 3'b101;
      // memory_array[29045] <= 3'b000;
      // memory_array[29046] <= 3'b111;
      // memory_array[29047] <= 3'b111;
      // memory_array[29048] <= 3'b111;
      // memory_array[29049] <= 3'b101;
      // memory_array[29050] <= 3'b101;
      // memory_array[29051] <= 3'b000;
      // memory_array[29052] <= 3'b111;
      // memory_array[29053] <= 3'b111;
      // memory_array[29054] <= 3'b101;
      // memory_array[29055] <= 3'b101;
      // memory_array[29056] <= 3'b000;
      // memory_array[29057] <= 3'b101;
      // memory_array[29058] <= 3'b101;
      // memory_array[29059] <= 3'b101;
      // memory_array[29060] <= 3'b000;
      // memory_array[29061] <= 3'b101;
      // memory_array[29062] <= 3'b000;
      // memory_array[29063] <= 3'b000;
      // memory_array[29064] <= 3'b101;
      // memory_array[29065] <= 3'b000;
      // memory_array[29066] <= 3'b111;
      // memory_array[29067] <= 3'b111;
      // memory_array[29068] <= 3'b111;
      // memory_array[29069] <= 3'b101;
      // memory_array[29070] <= 3'b000;
      // memory_array[29071] <= 3'b000;
      // memory_array[29072] <= 3'b101;
      // memory_array[29073] <= 3'b101;
      // memory_array[29074] <= 3'b101;
      // memory_array[29075] <= 3'b101;
      // memory_array[29076] <= 3'b101;
      // memory_array[29077] <= 3'b101;
      // memory_array[29078] <= 3'b000;
      // memory_array[29079] <= 3'b000;
      // memory_array[29080] <= 3'b000;
      // memory_array[29081] <= 3'b101;
      // memory_array[29082] <= 3'b000;
      // memory_array[29083] <= 3'b000;
      // memory_array[29084] <= 3'b101;
      // memory_array[29085] <= 3'b101;
      // memory_array[29086] <= 3'b000;
      // memory_array[29087] <= 3'b101;
      // memory_array[29088] <= 3'b101;
      // memory_array[29089] <= 3'b101;
      // memory_array[29090] <= 3'b101;
      // memory_array[29091] <= 3'b101;
      // memory_array[29092] <= 3'b101;
      // memory_array[29093] <= 3'b101;
      // memory_array[29094] <= 3'b101;
      // memory_array[29095] <= 3'b101;
      // memory_array[29096] <= 3'b101;
      // memory_array[29097] <= 3'b000;
      // memory_array[29098] <= 3'b101;
      // memory_array[29099] <= 3'b101;
      // memory_array[29100] <= 3'b000;
      // memory_array[29101] <= 3'b111;
      // memory_array[29102] <= 3'b101;
      // memory_array[29103] <= 3'b101;
      // memory_array[29104] <= 3'b101;
      // memory_array[29105] <= 3'b101;
      // memory_array[29106] <= 3'b101;
      // memory_array[29107] <= 3'b101;
      // memory_array[29108] <= 3'b101;
      // memory_array[29109] <= 3'b101;
      // memory_array[29110] <= 3'b101;
      // memory_array[29111] <= 3'b101;
      // memory_array[29112] <= 3'b000;
      // memory_array[29113] <= 3'b000;
      // memory_array[29114] <= 3'b101;
      // memory_array[29115] <= 3'b101;
      // memory_array[29116] <= 3'b101;
      // memory_array[29117] <= 3'b101;
      // memory_array[29118] <= 3'b101;
      // memory_array[29119] <= 3'b101;
      // memory_array[29120] <= 3'b000;
      // memory_array[29121] <= 3'b101;
      // memory_array[29122] <= 3'b101;
      // memory_array[29123] <= 3'b101;
      // memory_array[29124] <= 3'b101;
      // memory_array[29125] <= 3'b101;
      // memory_array[29126] <= 3'b101;
      // memory_array[29127] <= 3'b101;
      // memory_array[29128] <= 3'b101;
      // memory_array[29129] <= 3'b101;
      // memory_array[29130] <= 3'b101;
      // memory_array[29131] <= 3'b000;
      // memory_array[29132] <= 3'b101;
      // memory_array[29133] <= 3'b101;
      // memory_array[29134] <= 3'b101;
      // memory_array[29135] <= 3'b000;
      // memory_array[29136] <= 3'b101;
      // memory_array[29137] <= 3'b000;
      // memory_array[29138] <= 3'b000;
      // memory_array[29139] <= 3'b101;
      // memory_array[29140] <= 3'b000;
      // memory_array[29141] <= 3'b111;
      // memory_array[29142] <= 3'b101;
      // memory_array[29143] <= 3'b111;
      // memory_array[29144] <= 3'b101;
      // memory_array[29145] <= 3'b000;
      // memory_array[29146] <= 3'b000;
      // memory_array[29147] <= 3'b101;
      // memory_array[29148] <= 3'b101;
      // memory_array[29149] <= 3'b101;
      // memory_array[29150] <= 3'b101;
      // memory_array[29151] <= 3'b101;
      // memory_array[29152] <= 3'b101;
      // memory_array[29153] <= 3'b000;
      // memory_array[29154] <= 3'b000;
      // memory_array[29155] <= 3'b000;
      // memory_array[29156] <= 3'b101;
      // memory_array[29157] <= 3'b000;
      // memory_array[29158] <= 3'b000;
      // memory_array[29159] <= 3'b101;
      // memory_array[29160] <= 3'b101;
      // memory_array[29161] <= 3'b000;
      // memory_array[29162] <= 3'b101;
      // memory_array[29163] <= 3'b101;
      // memory_array[29164] <= 3'b101;
      // memory_array[29165] <= 3'b101;
      // memory_array[29166] <= 3'b101;
      // memory_array[29167] <= 3'b101;
      // memory_array[29168] <= 3'b101;
      // memory_array[29169] <= 3'b101;
      // memory_array[29170] <= 3'b101;
      // memory_array[29171] <= 3'b101;
      // memory_array[29172] <= 3'b000;
      // memory_array[29173] <= 3'b000;
      // memory_array[29174] <= 3'b101;
      // memory_array[29175] <= 3'b101;
      // memory_array[29176] <= 3'b000;
      // memory_array[29177] <= 3'b000;
      // memory_array[29178] <= 3'b000;
      // memory_array[29179] <= 3'b101;
      // memory_array[29180] <= 3'b000;
      // memory_array[29181] <= 3'b101;
      // memory_array[29182] <= 3'b000;
      // memory_array[29183] <= 3'b000;
      // memory_array[29184] <= 3'b101;
      // memory_array[29185] <= 3'b000;
      // memory_array[29186] <= 3'b111;
      // memory_array[29187] <= 3'b101;
      // memory_array[29188] <= 3'b111;
      // memory_array[29189] <= 3'b101;
      // memory_array[29190] <= 3'b101;
      // memory_array[29191] <= 3'b101;
      // memory_array[29192] <= 3'b111;
      // memory_array[29193] <= 3'b101;
      // memory_array[29194] <= 3'b101;
      // memory_array[29195] <= 3'b111;
      // memory_array[29196] <= 3'b111;
      // memory_array[29197] <= 3'b101;
      // memory_array[29198] <= 3'b101;
      // memory_array[29199] <= 3'b111;
      // memory_array[29200] <= 3'b111;
      // memory_array[29201] <= 3'b111;
      // memory_array[29202] <= 3'b111;
      // memory_array[29203] <= 3'b111;
      // memory_array[29204] <= 3'b101;
      // memory_array[29205] <= 3'b111;
      // memory_array[29206] <= 3'b111;
      // memory_array[29207] <= 3'b111;
      // memory_array[29208] <= 3'b101;
      // memory_array[29209] <= 3'b101;
      // memory_array[29210] <= 3'b101;
      // memory_array[29211] <= 3'b101;
      // memory_array[29212] <= 3'b101;
      // memory_array[29213] <= 3'b000;
      // memory_array[29214] <= 3'b101;
      // memory_array[29215] <= 3'b101;
      // memory_array[29216] <= 3'b000;
      // memory_array[29217] <= 3'b111;
      // memory_array[29218] <= 3'b101;
      // memory_array[29219] <= 3'b000;
      // memory_array[29220] <= 3'b000;
      // memory_array[29221] <= 3'b000;
      // memory_array[29222] <= 3'b101;
      // memory_array[29223] <= 3'b101;
      // memory_array[29224] <= 3'b101;
      // memory_array[29225] <= 3'b101;
      // memory_array[29226] <= 3'b000;
      // memory_array[29227] <= 3'b000;
      // memory_array[29228] <= 3'b000;
      // memory_array[29229] <= 3'b101;
      // memory_array[29230] <= 3'b101;
      // memory_array[29231] <= 3'b101;
      // memory_array[29232] <= 3'b101;
      // memory_array[29233] <= 3'b101;
      // memory_array[29234] <= 3'b101;
      // memory_array[29235] <= 3'b101;
      // memory_array[29236] <= 3'b101;
      // memory_array[29237] <= 3'b000;
      // memory_array[29238] <= 3'b101;
      // memory_array[29239] <= 3'b111;
      // memory_array[29240] <= 3'b101;
      // memory_array[29241] <= 3'b000;
      // memory_array[29242] <= 3'b101;
      // memory_array[29243] <= 3'b101;
      // memory_array[29244] <= 3'b101;
      // memory_array[29245] <= 3'b101;
      // memory_array[29246] <= 3'b101;
      // memory_array[29247] <= 3'b101;
      // memory_array[29248] <= 3'b101;
      // memory_array[29249] <= 3'b101;
      // memory_array[29250] <= 3'b101;
      // memory_array[29251] <= 3'b101;
      // memory_array[29252] <= 3'b000;
      // memory_array[29253] <= 3'b000;
      // memory_array[29254] <= 3'b101;
      // memory_array[29255] <= 3'b101;
      // memory_array[29256] <= 3'b101;
      // memory_array[29257] <= 3'b111;
      // memory_array[29258] <= 3'b000;
      // memory_array[29259] <= 3'b101;
      // memory_array[29260] <= 3'b101;
      // memory_array[29261] <= 3'b000;
      // memory_array[29262] <= 3'b111;
      // memory_array[29263] <= 3'b101;
      // memory_array[29264] <= 3'b000;
      // memory_array[29265] <= 3'b000;
      // memory_array[29266] <= 3'b000;
      // memory_array[29267] <= 3'b101;
      // memory_array[29268] <= 3'b101;
      // memory_array[29269] <= 3'b000;
      // memory_array[29270] <= 3'b101;
      // memory_array[29271] <= 3'b000;
      // memory_array[29272] <= 3'b101;
      // memory_array[29273] <= 3'b101;
      // memory_array[29274] <= 3'b101;
      // memory_array[29275] <= 3'b101;
      // memory_array[29276] <= 3'b101;
      // memory_array[29277] <= 3'b101;
      // memory_array[29278] <= 3'b101;
      // memory_array[29279] <= 3'b101;
      // memory_array[29280] <= 3'b101;
      // memory_array[29281] <= 3'b101;
      // memory_array[29282] <= 3'b000;
      // memory_array[29283] <= 3'b000;
      // memory_array[29284] <= 3'b000;
      // memory_array[29285] <= 3'b101;
      // memory_array[29286] <= 3'b000;
      // memory_array[29287] <= 3'b101;
      // memory_array[29288] <= 3'b101;
      // memory_array[29289] <= 3'b101;
      // memory_array[29290] <= 3'b101;
      // memory_array[29291] <= 3'b101;
      // memory_array[29292] <= 3'b101;
      // memory_array[29293] <= 3'b101;
      // memory_array[29294] <= 3'b101;
      // memory_array[29295] <= 3'b101;
      // memory_array[29296] <= 3'b000;
      // memory_array[29297] <= 3'b111;
      // memory_array[29298] <= 3'b101;
      // memory_array[29299] <= 3'b101;
      // memory_array[29300] <= 3'b101;
      // memory_array[29301] <= 3'b000;
      // memory_array[29302] <= 3'b000;
      // memory_array[29303] <= 3'b000;
      // memory_array[29304] <= 3'b101;
      // memory_array[29305] <= 3'b101;
      // memory_array[29306] <= 3'b101;
      // memory_array[29307] <= 3'b101;
      // memory_array[29308] <= 3'b101;
      // memory_array[29309] <= 3'b101;
      // memory_array[29310] <= 3'b101;
      // memory_array[29311] <= 3'b101;
      // memory_array[29312] <= 3'b000;
      // memory_array[29313] <= 3'b101;
      // memory_array[29314] <= 3'b111;
      // memory_array[29315] <= 3'b101;
      // memory_array[29316] <= 3'b000;
      // memory_array[29317] <= 3'b101;
      // memory_array[29318] <= 3'b101;
      // memory_array[29319] <= 3'b101;
      // memory_array[29320] <= 3'b101;
      // memory_array[29321] <= 3'b101;
      // memory_array[29322] <= 3'b101;
      // memory_array[29323] <= 3'b101;
      // memory_array[29324] <= 3'b101;
      // memory_array[29325] <= 3'b101;
      // memory_array[29326] <= 3'b101;
      // memory_array[29327] <= 3'b000;
      // memory_array[29328] <= 3'b000;
      // memory_array[29329] <= 3'b101;
      // memory_array[29330] <= 3'b101;
      // memory_array[29331] <= 3'b101;
      // memory_array[29332] <= 3'b111;
      // memory_array[29333] <= 3'b000;
      // memory_array[29334] <= 3'b101;
      // memory_array[29335] <= 3'b101;
      // memory_array[29336] <= 3'b000;
      // memory_array[29337] <= 3'b111;
      // memory_array[29338] <= 3'b101;
      // memory_array[29339] <= 3'b000;
      // memory_array[29340] <= 3'b000;
      // memory_array[29341] <= 3'b000;
      // memory_array[29342] <= 3'b101;
      // memory_array[29343] <= 3'b101;
      // memory_array[29344] <= 3'b000;
      // memory_array[29345] <= 3'b101;
      // memory_array[29346] <= 3'b000;
      // memory_array[29347] <= 3'b101;
      // memory_array[29348] <= 3'b101;
      // memory_array[29349] <= 3'b101;
      // memory_array[29350] <= 3'b101;
      // memory_array[29351] <= 3'b101;
      // memory_array[29352] <= 3'b101;
      // memory_array[29353] <= 3'b101;
      // memory_array[29354] <= 3'b101;
      // memory_array[29355] <= 3'b101;
      // memory_array[29356] <= 3'b101;
      // memory_array[29357] <= 3'b000;
      // memory_array[29358] <= 3'b000;
      // memory_array[29359] <= 3'b000;
      // memory_array[29360] <= 3'b101;
      // memory_array[29361] <= 3'b000;
      // memory_array[29362] <= 3'b101;
      // memory_array[29363] <= 3'b101;
      // memory_array[29364] <= 3'b101;
      // memory_array[29365] <= 3'b101;
      // memory_array[29366] <= 3'b101;
      // memory_array[29367] <= 3'b101;
      // memory_array[29368] <= 3'b101;
      // memory_array[29369] <= 3'b101;
      // memory_array[29370] <= 3'b101;
      // memory_array[29371] <= 3'b000;
      // memory_array[29372] <= 3'b111;
      // memory_array[29373] <= 3'b101;
      // memory_array[29374] <= 3'b101;
      // memory_array[29375] <= 3'b101;
      // memory_array[29376] <= 3'b101;
      // memory_array[29377] <= 3'b101;
      // memory_array[29378] <= 3'b000;
      // memory_array[29379] <= 3'b101;
      // memory_array[29380] <= 3'b101;
      // memory_array[29381] <= 3'b000;
      // memory_array[29382] <= 3'b111;
      // memory_array[29383] <= 3'b101;
      // memory_array[29384] <= 3'b000;
      // memory_array[29385] <= 3'b000;
      // memory_array[29386] <= 3'b000;
      // memory_array[29387] <= 3'b101;
      // memory_array[29388] <= 3'b101;
      // memory_array[29389] <= 3'b101;
      // memory_array[29390] <= 3'b101;
      // memory_array[29391] <= 3'b101;
      // memory_array[29392] <= 3'b111;
      // memory_array[29393] <= 3'b101;
      // memory_array[29394] <= 3'b101;
      // memory_array[29395] <= 3'b111;
      // memory_array[29396] <= 3'b111;
      // memory_array[29397] <= 3'b101;
      // memory_array[29398] <= 3'b101;
      // memory_array[29399] <= 3'b111;
      // memory_array[29400] <= 3'b111;
      // memory_array[29401] <= 3'b111;
      // memory_array[29402] <= 3'b111;
      // memory_array[29403] <= 3'b111;
      // memory_array[29404] <= 3'b111;
      // memory_array[29405] <= 3'b111;
      // memory_array[29406] <= 3'b111;
      // memory_array[29407] <= 3'b111;
      // memory_array[29408] <= 3'b101;
      // memory_array[29409] <= 3'b101;
      // memory_array[29410] <= 3'b101;
      // memory_array[29411] <= 3'b101;
      // memory_array[29412] <= 3'b000;
      // memory_array[29413] <= 3'b000;
      // memory_array[29414] <= 3'b000;
      // memory_array[29415] <= 3'b101;
      // memory_array[29416] <= 3'b000;
      // memory_array[29417] <= 3'b000;
      // memory_array[29418] <= 3'b000;
      // memory_array[29419] <= 3'b000;
      // memory_array[29420] <= 3'b101;
      // memory_array[29421] <= 3'b000;
      // memory_array[29422] <= 3'b101;
      // memory_array[29423] <= 3'b101;
      // memory_array[29424] <= 3'b101;
      // memory_array[29425] <= 3'b101;
      // memory_array[29426] <= 3'b000;
      // memory_array[29427] <= 3'b000;
      // memory_array[29428] <= 3'b000;
      // memory_array[29429] <= 3'b101;
      // memory_array[29430] <= 3'b000;
      // memory_array[29431] <= 3'b101;
      // memory_array[29432] <= 3'b000;
      // memory_array[29433] <= 3'b000;
      // memory_array[29434] <= 3'b000;
      // memory_array[29435] <= 3'b101;
      // memory_array[29436] <= 3'b101;
      // memory_array[29437] <= 3'b101;
      // memory_array[29438] <= 3'b101;
      // memory_array[29439] <= 3'b000;
      // memory_array[29440] <= 3'b000;
      // memory_array[29441] <= 3'b101;
      // memory_array[29442] <= 3'b000;
      // memory_array[29443] <= 3'b000;
      // memory_array[29444] <= 3'b101;
      // memory_array[29445] <= 3'b101;
      // memory_array[29446] <= 3'b101;
      // memory_array[29447] <= 3'b101;
      // memory_array[29448] <= 3'b101;
      // memory_array[29449] <= 3'b101;
      // memory_array[29450] <= 3'b101;
      // memory_array[29451] <= 3'b101;
      // memory_array[29452] <= 3'b101;
      // memory_array[29453] <= 3'b101;
      // memory_array[29454] <= 3'b000;
      // memory_array[29455] <= 3'b000;
      // memory_array[29456] <= 3'b101;
      // memory_array[29457] <= 3'b000;
      // memory_array[29458] <= 3'b101;
      // memory_array[29459] <= 3'b101;
      // memory_array[29460] <= 3'b101;
      // memory_array[29461] <= 3'b000;
      // memory_array[29462] <= 3'b000;
      // memory_array[29463] <= 3'b000;
      // memory_array[29464] <= 3'b000;
      // memory_array[29465] <= 3'b101;
      // memory_array[29466] <= 3'b000;
      // memory_array[29467] <= 3'b101;
      // memory_array[29468] <= 3'b000;
      // memory_array[29469] <= 3'b101;
      // memory_array[29470] <= 3'b000;
      // memory_array[29471] <= 3'b101;
      // memory_array[29472] <= 3'b101;
      // memory_array[29473] <= 3'b000;
      // memory_array[29474] <= 3'b101;
      // memory_array[29475] <= 3'b101;
      // memory_array[29476] <= 3'b101;
      // memory_array[29477] <= 3'b101;
      // memory_array[29478] <= 3'b101;
      // memory_array[29479] <= 3'b101;
      // memory_array[29480] <= 3'b101;
      // memory_array[29481] <= 3'b000;
      // memory_array[29482] <= 3'b101;
      // memory_array[29483] <= 3'b101;
      // memory_array[29484] <= 3'b000;
      // memory_array[29485] <= 3'b000;
      // memory_array[29486] <= 3'b000;
      // memory_array[29487] <= 3'b000;
      // memory_array[29488] <= 3'b000;
      // memory_array[29489] <= 3'b101;
      // memory_array[29490] <= 3'b000;
      // memory_array[29491] <= 3'b101;
      // memory_array[29492] <= 3'b000;
      // memory_array[29493] <= 3'b000;
      // memory_array[29494] <= 3'b000;
      // memory_array[29495] <= 3'b101;
      // memory_array[29496] <= 3'b101;
      // memory_array[29497] <= 3'b101;
      // memory_array[29498] <= 3'b101;
      // memory_array[29499] <= 3'b101;
      // memory_array[29500] <= 3'b101;
      // memory_array[29501] <= 3'b000;
      // memory_array[29502] <= 3'b000;
      // memory_array[29503] <= 3'b000;
      // memory_array[29504] <= 3'b101;
      // memory_array[29505] <= 3'b000;
      // memory_array[29506] <= 3'b101;
      // memory_array[29507] <= 3'b000;
      // memory_array[29508] <= 3'b000;
      // memory_array[29509] <= 3'b000;
      // memory_array[29510] <= 3'b101;
      // memory_array[29511] <= 3'b101;
      // memory_array[29512] <= 3'b101;
      // memory_array[29513] <= 3'b101;
      // memory_array[29514] <= 3'b000;
      // memory_array[29515] <= 3'b000;
      // memory_array[29516] <= 3'b101;
      // memory_array[29517] <= 3'b000;
      // memory_array[29518] <= 3'b000;
      // memory_array[29519] <= 3'b101;
      // memory_array[29520] <= 3'b101;
      // memory_array[29521] <= 3'b101;
      // memory_array[29522] <= 3'b101;
      // memory_array[29523] <= 3'b101;
      // memory_array[29524] <= 3'b101;
      // memory_array[29525] <= 3'b101;
      // memory_array[29526] <= 3'b101;
      // memory_array[29527] <= 3'b101;
      // memory_array[29528] <= 3'b101;
      // memory_array[29529] <= 3'b000;
      // memory_array[29530] <= 3'b000;
      // memory_array[29531] <= 3'b101;
      // memory_array[29532] <= 3'b000;
      // memory_array[29533] <= 3'b101;
      // memory_array[29534] <= 3'b101;
      // memory_array[29535] <= 3'b101;
      // memory_array[29536] <= 3'b000;
      // memory_array[29537] <= 3'b000;
      // memory_array[29538] <= 3'b000;
      // memory_array[29539] <= 3'b000;
      // memory_array[29540] <= 3'b101;
      // memory_array[29541] <= 3'b000;
      // memory_array[29542] <= 3'b101;
      // memory_array[29543] <= 3'b000;
      // memory_array[29544] <= 3'b101;
      // memory_array[29545] <= 3'b000;
      // memory_array[29546] <= 3'b101;
      // memory_array[29547] <= 3'b101;
      // memory_array[29548] <= 3'b000;
      // memory_array[29549] <= 3'b101;
      // memory_array[29550] <= 3'b101;
      // memory_array[29551] <= 3'b101;
      // memory_array[29552] <= 3'b101;
      // memory_array[29553] <= 3'b101;
      // memory_array[29554] <= 3'b101;
      // memory_array[29555] <= 3'b101;
      // memory_array[29556] <= 3'b000;
      // memory_array[29557] <= 3'b101;
      // memory_array[29558] <= 3'b101;
      // memory_array[29559] <= 3'b000;
      // memory_array[29560] <= 3'b000;
      // memory_array[29561] <= 3'b000;
      // memory_array[29562] <= 3'b000;
      // memory_array[29563] <= 3'b000;
      // memory_array[29564] <= 3'b101;
      // memory_array[29565] <= 3'b000;
      // memory_array[29566] <= 3'b101;
      // memory_array[29567] <= 3'b000;
      // memory_array[29568] <= 3'b000;
      // memory_array[29569] <= 3'b000;
      // memory_array[29570] <= 3'b101;
      // memory_array[29571] <= 3'b101;
      // memory_array[29572] <= 3'b101;
      // memory_array[29573] <= 3'b101;
      // memory_array[29574] <= 3'b101;
      // memory_array[29575] <= 3'b101;
      // memory_array[29576] <= 3'b101;
      // memory_array[29577] <= 3'b000;
      // memory_array[29578] <= 3'b000;
      // memory_array[29579] <= 3'b000;
      // memory_array[29580] <= 3'b101;
      // memory_array[29581] <= 3'b000;
      // memory_array[29582] <= 3'b000;
      // memory_array[29583] <= 3'b000;
      // memory_array[29584] <= 3'b000;
      // memory_array[29585] <= 3'b101;
      // memory_array[29586] <= 3'b000;
      // memory_array[29587] <= 3'b101;
      // memory_array[29588] <= 3'b101;
      // memory_array[29589] <= 3'b101;
      // memory_array[29590] <= 3'b101;
      // memory_array[29591] <= 3'b101;
      // memory_array[29592] <= 3'b111;
      // memory_array[29593] <= 3'b111;
      // memory_array[29594] <= 3'b111;
      // memory_array[29595] <= 3'b101;
      // memory_array[29596] <= 3'b101;
      // memory_array[29597] <= 3'b111;
      // memory_array[29598] <= 3'b111;
      // memory_array[29599] <= 3'b111;
      // memory_array[29600] <= 3'b111;
      // memory_array[29601] <= 3'b111;
      // memory_array[29602] <= 3'b111;
      // memory_array[29603] <= 3'b101;
      // memory_array[29604] <= 3'b111;
      // memory_array[29605] <= 3'b111;
      // memory_array[29606] <= 3'b111;
      // memory_array[29607] <= 3'b111;
      // memory_array[29608] <= 3'b101;
      // memory_array[29609] <= 3'b101;
      // memory_array[29610] <= 3'b101;
      // memory_array[29611] <= 3'b101;
      // memory_array[29612] <= 3'b000;
      // memory_array[29613] <= 3'b000;
      // memory_array[29614] <= 3'b000;
      // memory_array[29615] <= 3'b000;
      // memory_array[29616] <= 3'b101;
      // memory_array[29617] <= 3'b101;
      // memory_array[29618] <= 3'b000;
      // memory_array[29619] <= 3'b111;
      // memory_array[29620] <= 3'b000;
      // memory_array[29621] <= 3'b111;
      // memory_array[29622] <= 3'b101;
      // memory_array[29623] <= 3'b101;
      // memory_array[29624] <= 3'b101;
      // memory_array[29625] <= 3'b101;
      // memory_array[29626] <= 3'b101;
      // memory_array[29627] <= 3'b000;
      // memory_array[29628] <= 3'b000;
      // memory_array[29629] <= 3'b000;
      // memory_array[29630] <= 3'b000;
      // memory_array[29631] <= 3'b101;
      // memory_array[29632] <= 3'b101;
      // memory_array[29633] <= 3'b000;
      // memory_array[29634] <= 3'b000;
      // memory_array[29635] <= 3'b000;
      // memory_array[29636] <= 3'b000;
      // memory_array[29637] <= 3'b000;
      // memory_array[29638] <= 3'b000;
      // memory_array[29639] <= 3'b101;
      // memory_array[29640] <= 3'b101;
      // memory_array[29641] <= 3'b101;
      // memory_array[29642] <= 3'b000;
      // memory_array[29643] <= 3'b000;
      // memory_array[29644] <= 3'b000;
      // memory_array[29645] <= 3'b000;
      // memory_array[29646] <= 3'b000;
      // memory_array[29647] <= 3'b000;
      // memory_array[29648] <= 3'b000;
      // memory_array[29649] <= 3'b000;
      // memory_array[29650] <= 3'b000;
      // memory_array[29651] <= 3'b000;
      // memory_array[29652] <= 3'b000;
      // memory_array[29653] <= 3'b000;
      // memory_array[29654] <= 3'b000;
      // memory_array[29655] <= 3'b000;
      // memory_array[29656] <= 3'b000;
      // memory_array[29657] <= 3'b000;
      // memory_array[29658] <= 3'b000;
      // memory_array[29659] <= 3'b000;
      // memory_array[29660] <= 3'b000;
      // memory_array[29661] <= 3'b101;
      // memory_array[29662] <= 3'b101;
      // memory_array[29663] <= 3'b000;
      // memory_array[29664] <= 3'b111;
      // memory_array[29665] <= 3'b000;
      // memory_array[29666] <= 3'b101;
      // memory_array[29667] <= 3'b101;
      // memory_array[29668] <= 3'b000;
      // memory_array[29669] <= 3'b000;
      // memory_array[29670] <= 3'b000;
      // memory_array[29671] <= 3'b000;
      // memory_array[29672] <= 3'b000;
      // memory_array[29673] <= 3'b000;
      // memory_array[29674] <= 3'b000;
      // memory_array[29675] <= 3'b000;
      // memory_array[29676] <= 3'b000;
      // memory_array[29677] <= 3'b000;
      // memory_array[29678] <= 3'b000;
      // memory_array[29679] <= 3'b000;
      // memory_array[29680] <= 3'b000;
      // memory_array[29681] <= 3'b000;
      // memory_array[29682] <= 3'b101;
      // memory_array[29683] <= 3'b101;
      // memory_array[29684] <= 3'b101;
      // memory_array[29685] <= 3'b101;
      // memory_array[29686] <= 3'b000;
      // memory_array[29687] <= 3'b000;
      // memory_array[29688] <= 3'b000;
      // memory_array[29689] <= 3'b000;
      // memory_array[29690] <= 3'b000;
      // memory_array[29691] <= 3'b101;
      // memory_array[29692] <= 3'b101;
      // memory_array[29693] <= 3'b000;
      // memory_array[29694] <= 3'b000;
      // memory_array[29695] <= 3'b000;
      // memory_array[29696] <= 3'b000;
      // memory_array[29697] <= 3'b101;
      // memory_array[29698] <= 3'b101;
      // memory_array[29699] <= 3'b101;
      // memory_array[29700] <= 3'b101;
      // memory_array[29701] <= 3'b101;
      // memory_array[29702] <= 3'b000;
      // memory_array[29703] <= 3'b000;
      // memory_array[29704] <= 3'b000;
      // memory_array[29705] <= 3'b000;
      // memory_array[29706] <= 3'b101;
      // memory_array[29707] <= 3'b101;
      // memory_array[29708] <= 3'b000;
      // memory_array[29709] <= 3'b000;
      // memory_array[29710] <= 3'b000;
      // memory_array[29711] <= 3'b000;
      // memory_array[29712] <= 3'b000;
      // memory_array[29713] <= 3'b000;
      // memory_array[29714] <= 3'b101;
      // memory_array[29715] <= 3'b101;
      // memory_array[29716] <= 3'b101;
      // memory_array[29717] <= 3'b000;
      // memory_array[29718] <= 3'b000;
      // memory_array[29719] <= 3'b000;
      // memory_array[29720] <= 3'b000;
      // memory_array[29721] <= 3'b000;
      // memory_array[29722] <= 3'b000;
      // memory_array[29723] <= 3'b000;
      // memory_array[29724] <= 3'b000;
      // memory_array[29725] <= 3'b000;
      // memory_array[29726] <= 3'b000;
      // memory_array[29727] <= 3'b000;
      // memory_array[29728] <= 3'b000;
      // memory_array[29729] <= 3'b000;
      // memory_array[29730] <= 3'b000;
      // memory_array[29731] <= 3'b000;
      // memory_array[29732] <= 3'b000;
      // memory_array[29733] <= 3'b000;
      // memory_array[29734] <= 3'b000;
      // memory_array[29735] <= 3'b000;
      // memory_array[29736] <= 3'b101;
      // memory_array[29737] <= 3'b101;
      // memory_array[29738] <= 3'b000;
      // memory_array[29739] <= 3'b111;
      // memory_array[29740] <= 3'b000;
      // memory_array[29741] <= 3'b101;
      // memory_array[29742] <= 3'b101;
      // memory_array[29743] <= 3'b000;
      // memory_array[29744] <= 3'b000;
      // memory_array[29745] <= 3'b000;
      // memory_array[29746] <= 3'b000;
      // memory_array[29747] <= 3'b000;
      // memory_array[29748] <= 3'b000;
      // memory_array[29749] <= 3'b000;
      // memory_array[29750] <= 3'b000;
      // memory_array[29751] <= 3'b000;
      // memory_array[29752] <= 3'b000;
      // memory_array[29753] <= 3'b000;
      // memory_array[29754] <= 3'b000;
      // memory_array[29755] <= 3'b000;
      // memory_array[29756] <= 3'b000;
      // memory_array[29757] <= 3'b101;
      // memory_array[29758] <= 3'b101;
      // memory_array[29759] <= 3'b101;
      // memory_array[29760] <= 3'b101;
      // memory_array[29761] <= 3'b000;
      // memory_array[29762] <= 3'b000;
      // memory_array[29763] <= 3'b000;
      // memory_array[29764] <= 3'b000;
      // memory_array[29765] <= 3'b000;
      // memory_array[29766] <= 3'b101;
      // memory_array[29767] <= 3'b101;
      // memory_array[29768] <= 3'b000;
      // memory_array[29769] <= 3'b000;
      // memory_array[29770] <= 3'b000;
      // memory_array[29771] <= 3'b000;
      // memory_array[29772] <= 3'b101;
      // memory_array[29773] <= 3'b101;
      // memory_array[29774] <= 3'b101;
      // memory_array[29775] <= 3'b101;
      // memory_array[29776] <= 3'b101;
      // memory_array[29777] <= 3'b000;
      // memory_array[29778] <= 3'b000;
      // memory_array[29779] <= 3'b000;
      // memory_array[29780] <= 3'b000;
      // memory_array[29781] <= 3'b101;
      // memory_array[29782] <= 3'b101;
      // memory_array[29783] <= 3'b000;
      // memory_array[29784] <= 3'b111;
      // memory_array[29785] <= 3'b000;
      // memory_array[29786] <= 3'b111;
      // memory_array[29787] <= 3'b101;
      // memory_array[29788] <= 3'b101;
      // memory_array[29789] <= 3'b101;
      // memory_array[29790] <= 3'b101;
      // memory_array[29791] <= 3'b101;
      // memory_array[29792] <= 3'b111;
      // memory_array[29793] <= 3'b111;
      // memory_array[29794] <= 3'b111;
      // memory_array[29795] <= 3'b101;
      // memory_array[29796] <= 3'b101;
      // memory_array[29797] <= 3'b111;
      // memory_array[29798] <= 3'b111;
      // memory_array[29799] <= 3'b111;
      // memory_array[29800] <= 3'b111;
      // memory_array[29801] <= 3'b111;
      // memory_array[29802] <= 3'b111;
      // memory_array[29803] <= 3'b111;
      // memory_array[29804] <= 3'b111;
      // memory_array[29805] <= 3'b111;
      // memory_array[29806] <= 3'b111;
      // memory_array[29807] <= 3'b111;
      // memory_array[29808] <= 3'b101;
      // memory_array[29809] <= 3'b101;
      // memory_array[29810] <= 3'b101;
      // memory_array[29811] <= 3'b101;
      // memory_array[29812] <= 3'b101;
      // memory_array[29813] <= 3'b101;
      // memory_array[29814] <= 3'b000;
      // memory_array[29815] <= 3'b101;
      // memory_array[29816] <= 3'b000;
      // memory_array[29817] <= 3'b000;
      // memory_array[29818] <= 3'b000;
      // memory_array[29819] <= 3'b000;
      // memory_array[29820] <= 3'b000;
      // memory_array[29821] <= 3'b101;
      // memory_array[29822] <= 3'b101;
      // memory_array[29823] <= 3'b101;
      // memory_array[29824] <= 3'b101;
      // memory_array[29825] <= 3'b101;
      // memory_array[29826] <= 3'b101;
      // memory_array[29827] <= 3'b101;
      // memory_array[29828] <= 3'b101;
      // memory_array[29829] <= 3'b101;
      // memory_array[29830] <= 3'b101;
      // memory_array[29831] <= 3'b101;
      // memory_array[29832] <= 3'b101;
      // memory_array[29833] <= 3'b101;
      // memory_array[29834] <= 3'b101;
      // memory_array[29835] <= 3'b101;
      // memory_array[29836] <= 3'b101;
      // memory_array[29837] <= 3'b101;
      // memory_array[29838] <= 3'b101;
      // memory_array[29839] <= 3'b101;
      // memory_array[29840] <= 3'b101;
      // memory_array[29841] <= 3'b101;
      // memory_array[29842] <= 3'b101;
      // memory_array[29843] <= 3'b101;
      // memory_array[29844] <= 3'b101;
      // memory_array[29845] <= 3'b101;
      // memory_array[29846] <= 3'b101;
      // memory_array[29847] <= 3'b101;
      // memory_array[29848] <= 3'b101;
      // memory_array[29849] <= 3'b101;
      // memory_array[29850] <= 3'b101;
      // memory_array[29851] <= 3'b101;
      // memory_array[29852] <= 3'b101;
      // memory_array[29853] <= 3'b101;
      // memory_array[29854] <= 3'b101;
      // memory_array[29855] <= 3'b101;
      // memory_array[29856] <= 3'b101;
      // memory_array[29857] <= 3'b101;
      // memory_array[29858] <= 3'b101;
      // memory_array[29859] <= 3'b000;
      // memory_array[29860] <= 3'b101;
      // memory_array[29861] <= 3'b000;
      // memory_array[29862] <= 3'b000;
      // memory_array[29863] <= 3'b000;
      // memory_array[29864] <= 3'b000;
      // memory_array[29865] <= 3'b000;
      // memory_array[29866] <= 3'b101;
      // memory_array[29867] <= 3'b101;
      // memory_array[29868] <= 3'b101;
      // memory_array[29869] <= 3'b101;
      // memory_array[29870] <= 3'b101;
      // memory_array[29871] <= 3'b101;
      // memory_array[29872] <= 3'b101;
      // memory_array[29873] <= 3'b101;
      // memory_array[29874] <= 3'b101;
      // memory_array[29875] <= 3'b101;
      // memory_array[29876] <= 3'b101;
      // memory_array[29877] <= 3'b101;
      // memory_array[29878] <= 3'b101;
      // memory_array[29879] <= 3'b101;
      // memory_array[29880] <= 3'b101;
      // memory_array[29881] <= 3'b101;
      // memory_array[29882] <= 3'b101;
      // memory_array[29883] <= 3'b101;
      // memory_array[29884] <= 3'b101;
      // memory_array[29885] <= 3'b101;
      // memory_array[29886] <= 3'b101;
      // memory_array[29887] <= 3'b101;
      // memory_array[29888] <= 3'b101;
      // memory_array[29889] <= 3'b101;
      // memory_array[29890] <= 3'b101;
      // memory_array[29891] <= 3'b101;
      // memory_array[29892] <= 3'b101;
      // memory_array[29893] <= 3'b101;
      // memory_array[29894] <= 3'b101;
      // memory_array[29895] <= 3'b101;
      // memory_array[29896] <= 3'b101;
      // memory_array[29897] <= 3'b101;
      // memory_array[29898] <= 3'b101;
      // memory_array[29899] <= 3'b101;
      // memory_array[29900] <= 3'b101;
      // memory_array[29901] <= 3'b101;
      // memory_array[29902] <= 3'b101;
      // memory_array[29903] <= 3'b101;
      // memory_array[29904] <= 3'b101;
      // memory_array[29905] <= 3'b101;
      // memory_array[29906] <= 3'b101;
      // memory_array[29907] <= 3'b101;
      // memory_array[29908] <= 3'b101;
      // memory_array[29909] <= 3'b101;
      // memory_array[29910] <= 3'b101;
      // memory_array[29911] <= 3'b101;
      // memory_array[29912] <= 3'b101;
      // memory_array[29913] <= 3'b101;
      // memory_array[29914] <= 3'b101;
      // memory_array[29915] <= 3'b101;
      // memory_array[29916] <= 3'b101;
      // memory_array[29917] <= 3'b101;
      // memory_array[29918] <= 3'b101;
      // memory_array[29919] <= 3'b101;
      // memory_array[29920] <= 3'b101;
      // memory_array[29921] <= 3'b101;
      // memory_array[29922] <= 3'b101;
      // memory_array[29923] <= 3'b101;
      // memory_array[29924] <= 3'b101;
      // memory_array[29925] <= 3'b101;
      // memory_array[29926] <= 3'b101;
      // memory_array[29927] <= 3'b101;
      // memory_array[29928] <= 3'b101;
      // memory_array[29929] <= 3'b101;
      // memory_array[29930] <= 3'b101;
      // memory_array[29931] <= 3'b101;
      // memory_array[29932] <= 3'b101;
      // memory_array[29933] <= 3'b101;
      // memory_array[29934] <= 3'b000;
      // memory_array[29935] <= 3'b101;
      // memory_array[29936] <= 3'b000;
      // memory_array[29937] <= 3'b000;
      // memory_array[29938] <= 3'b000;
      // memory_array[29939] <= 3'b000;
      // memory_array[29940] <= 3'b000;
      // memory_array[29941] <= 3'b101;
      // memory_array[29942] <= 3'b101;
      // memory_array[29943] <= 3'b101;
      // memory_array[29944] <= 3'b101;
      // memory_array[29945] <= 3'b101;
      // memory_array[29946] <= 3'b101;
      // memory_array[29947] <= 3'b101;
      // memory_array[29948] <= 3'b101;
      // memory_array[29949] <= 3'b101;
      // memory_array[29950] <= 3'b101;
      // memory_array[29951] <= 3'b101;
      // memory_array[29952] <= 3'b101;
      // memory_array[29953] <= 3'b101;
      // memory_array[29954] <= 3'b101;
      // memory_array[29955] <= 3'b101;
      // memory_array[29956] <= 3'b101;
      // memory_array[29957] <= 3'b101;
      // memory_array[29958] <= 3'b101;
      // memory_array[29959] <= 3'b101;
      // memory_array[29960] <= 3'b101;
      // memory_array[29961] <= 3'b101;
      // memory_array[29962] <= 3'b101;
      // memory_array[29963] <= 3'b101;
      // memory_array[29964] <= 3'b101;
      // memory_array[29965] <= 3'b101;
      // memory_array[29966] <= 3'b101;
      // memory_array[29967] <= 3'b101;
      // memory_array[29968] <= 3'b101;
      // memory_array[29969] <= 3'b101;
      // memory_array[29970] <= 3'b101;
      // memory_array[29971] <= 3'b101;
      // memory_array[29972] <= 3'b101;
      // memory_array[29973] <= 3'b101;
      // memory_array[29974] <= 3'b101;
      // memory_array[29975] <= 3'b101;
      // memory_array[29976] <= 3'b101;
      // memory_array[29977] <= 3'b101;
      // memory_array[29978] <= 3'b101;
      // memory_array[29979] <= 3'b000;
      // memory_array[29980] <= 3'b101;
      // memory_array[29981] <= 3'b000;
      // memory_array[29982] <= 3'b000;
      // memory_array[29983] <= 3'b000;
      // memory_array[29984] <= 3'b000;
      // memory_array[29985] <= 3'b000;
      // memory_array[29986] <= 3'b101;
      // memory_array[29987] <= 3'b101;
      // memory_array[29988] <= 3'b101;
      // memory_array[29989] <= 3'b101;
      // memory_array[29990] <= 3'b101;
      // memory_array[29991] <= 3'b101;
      // memory_array[29992] <= 3'b111;
      // memory_array[29993] <= 3'b111;
      // memory_array[29994] <= 3'b111;
      // memory_array[29995] <= 3'b111;
      // memory_array[29996] <= 3'b111;
      // memory_array[29997] <= 3'b111;
      // memory_array[29998] <= 3'b111;
      // memory_array[29999] <= 3'b111;

    end

    // <= : every line executed in parallel in always block
    always @(posedge clk_10mhz) begin
        // Display pixel.
        if (h_counter > 199)  // Horizontal blanking.
      	begin
      	  red <= 0;
          green <= 0;
          blue <= 0;
      	end else if (v_counter > 599)  // Vertical blanking.
      	begin
      	  red <= 0;
          green <= 0;
          blue <= 0;
      	end else // Active video.
        begin
          red <= memory_array[h_counter + ((v_counter / 4) * 200)][0];
          green <= memory_array[h_counter + ((v_counter / 4) * 200)][1];
          blue <= memory_array[h_counter + ((v_counter / 4) * 200)][2];
        end

        // Horitonal sync.
        if (h_counter > 209 && h_counter < 242)
        begin
          h_sync <= 1;
        end else
        begin
          h_sync <= 0;
        end

        // Vertical sync.
        if (v_counter > 600 && v_counter < 605)
        begin
          v_sync <= 1;
        end else
        begin
          v_sync <= 0;
        end

        // Increment / reset counters.
        h_counter <= h_counter + 1'b1;

        if (h_counter == 264)
        begin
          h_counter <= 0;
          v_counter <= v_counter + 1'b1;
        end

        if (v_counter == 628)
        begin
          v_counter <= 0;
        end
    end

endmodule
